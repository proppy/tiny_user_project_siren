magic
tech gf180mcuC
magscale 1 10
timestamp 1668865357
<< metal1 >>
rect 11890 47854 11902 47906
rect 11954 47903 11966 47906
rect 12786 47903 12798 47906
rect 11954 47857 12798 47903
rect 11954 47854 11966 47857
rect 12786 47854 12798 47857
rect 12850 47854 12862 47906
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 32398 46002 32450 46014
rect 42478 46002 42530 46014
rect 4050 45950 4062 46002
rect 4114 45950 4126 46002
rect 5954 45950 5966 46002
rect 6018 45950 6030 46002
rect 12786 45950 12798 46002
rect 12850 45950 12862 46002
rect 24434 45950 24446 46002
rect 24498 45950 24510 46002
rect 25330 45950 25342 46002
rect 25394 45950 25406 46002
rect 27458 45950 27470 46002
rect 27522 45950 27534 46002
rect 33842 45950 33854 46002
rect 33906 45950 33918 46002
rect 35746 45950 35758 46002
rect 35810 45950 35822 46002
rect 43698 45950 43710 46002
rect 43762 45950 43774 46002
rect 32398 45938 32450 45950
rect 42478 45938 42530 45950
rect 31950 45890 32002 45902
rect 4946 45838 4958 45890
rect 5010 45838 5022 45890
rect 8754 45838 8766 45890
rect 8818 45838 8830 45890
rect 9986 45838 9998 45890
rect 10050 45838 10062 45890
rect 13570 45838 13582 45890
rect 13634 45838 13646 45890
rect 15922 45838 15934 45890
rect 15986 45838 15998 45890
rect 16482 45838 16494 45890
rect 16546 45838 16558 45890
rect 19954 45838 19966 45890
rect 20018 45838 20030 45890
rect 20626 45838 20638 45890
rect 20690 45838 20702 45890
rect 21298 45838 21310 45890
rect 21362 45838 21374 45890
rect 22082 45838 22094 45890
rect 22146 45838 22158 45890
rect 28242 45838 28254 45890
rect 28306 45838 28318 45890
rect 31378 45838 31390 45890
rect 31442 45838 31454 45890
rect 33170 45838 33182 45890
rect 33234 45838 33246 45890
rect 35074 45838 35086 45890
rect 35138 45838 35150 45890
rect 42914 45838 42926 45890
rect 42978 45838 42990 45890
rect 31950 45826 32002 45838
rect 2270 45778 2322 45790
rect 2270 45714 2322 45726
rect 2942 45778 2994 45790
rect 29262 45778 29314 45790
rect 8082 45726 8094 45778
rect 8146 45726 8158 45778
rect 10658 45726 10670 45778
rect 10722 45726 10734 45778
rect 2942 45714 2994 45726
rect 29262 45714 29314 45726
rect 29486 45778 29538 45790
rect 29486 45714 29538 45726
rect 29822 45778 29874 45790
rect 29822 45714 29874 45726
rect 30382 45778 30434 45790
rect 30382 45714 30434 45726
rect 31166 45778 31218 45790
rect 31166 45714 31218 45726
rect 37886 45778 37938 45790
rect 37886 45714 37938 45726
rect 39902 45778 39954 45790
rect 39902 45714 39954 45726
rect 48078 45778 48130 45790
rect 48078 45714 48130 45726
rect 1822 45666 1874 45678
rect 29598 45666 29650 45678
rect 17490 45614 17502 45666
rect 17554 45614 17566 45666
rect 1822 45602 1874 45614
rect 29598 45602 29650 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 1822 45330 1874 45342
rect 1822 45266 1874 45278
rect 2494 45330 2546 45342
rect 2494 45266 2546 45278
rect 3166 45330 3218 45342
rect 3166 45266 3218 45278
rect 3502 45330 3554 45342
rect 3502 45266 3554 45278
rect 5518 45330 5570 45342
rect 24446 45330 24498 45342
rect 12226 45278 12238 45330
rect 12290 45278 12302 45330
rect 23762 45278 23774 45330
rect 23826 45278 23838 45330
rect 5518 45266 5570 45278
rect 24446 45266 24498 45278
rect 26238 45330 26290 45342
rect 26238 45266 26290 45278
rect 27022 45330 27074 45342
rect 27022 45266 27074 45278
rect 30718 45330 30770 45342
rect 30718 45266 30770 45278
rect 31166 45330 31218 45342
rect 31166 45266 31218 45278
rect 33518 45330 33570 45342
rect 33518 45266 33570 45278
rect 34750 45330 34802 45342
rect 34750 45266 34802 45278
rect 18398 45218 18450 45230
rect 6850 45166 6862 45218
rect 6914 45166 6926 45218
rect 18398 45154 18450 45166
rect 27134 45218 27186 45230
rect 27134 45154 27186 45166
rect 27358 45218 27410 45230
rect 27358 45154 27410 45166
rect 29150 45218 29202 45230
rect 29150 45154 29202 45166
rect 29374 45218 29426 45230
rect 29374 45154 29426 45166
rect 30046 45218 30098 45230
rect 30046 45154 30098 45166
rect 30606 45218 30658 45230
rect 30606 45154 30658 45166
rect 31614 45218 31666 45230
rect 31614 45154 31666 45166
rect 10110 45106 10162 45118
rect 6178 45054 6190 45106
rect 6242 45054 6254 45106
rect 9762 45054 9774 45106
rect 9826 45054 9838 45106
rect 10110 45042 10162 45054
rect 10334 45106 10386 45118
rect 10334 45042 10386 45054
rect 11006 45106 11058 45118
rect 11006 45042 11058 45054
rect 11118 45106 11170 45118
rect 11118 45042 11170 45054
rect 11230 45106 11282 45118
rect 17726 45106 17778 45118
rect 14578 45054 14590 45106
rect 14642 45054 14654 45106
rect 15362 45054 15374 45106
rect 15426 45054 15438 45106
rect 16370 45054 16382 45106
rect 16434 45054 16446 45106
rect 11230 45042 11282 45054
rect 17726 45042 17778 45054
rect 17950 45106 18002 45118
rect 17950 45042 18002 45054
rect 18174 45106 18226 45118
rect 24222 45106 24274 45118
rect 18946 45054 18958 45106
rect 19010 45054 19022 45106
rect 20850 45054 20862 45106
rect 20914 45054 20926 45106
rect 21410 45054 21422 45106
rect 21474 45054 21486 45106
rect 18174 45042 18226 45054
rect 24222 45042 24274 45054
rect 24558 45106 24610 45118
rect 24558 45042 24610 45054
rect 24782 45106 24834 45118
rect 24782 45042 24834 45054
rect 25566 45106 25618 45118
rect 25566 45042 25618 45054
rect 26014 45106 26066 45118
rect 26014 45042 26066 45054
rect 26126 45106 26178 45118
rect 26126 45042 26178 45054
rect 26686 45106 26738 45118
rect 26686 45042 26738 45054
rect 27918 45106 27970 45118
rect 27918 45042 27970 45054
rect 28142 45106 28194 45118
rect 32510 45106 32562 45118
rect 28466 45054 28478 45106
rect 28530 45054 28542 45106
rect 28142 45042 28194 45054
rect 32510 45042 32562 45054
rect 4062 44994 4114 45006
rect 4062 44930 4114 44942
rect 4510 44994 4562 45006
rect 4510 44930 4562 44942
rect 4958 44994 5010 45006
rect 4958 44930 5010 44942
rect 5406 44994 5458 45006
rect 10222 44994 10274 45006
rect 8978 44942 8990 44994
rect 9042 44942 9054 44994
rect 5406 44930 5458 44942
rect 10222 44930 10274 44942
rect 11454 44994 11506 45006
rect 11454 44930 11506 44942
rect 15934 44994 15986 45006
rect 28030 44994 28082 45006
rect 29934 44994 29986 45006
rect 16258 44942 16270 44994
rect 16322 44942 16334 44994
rect 19954 44942 19966 44994
rect 20018 44942 20030 44994
rect 29026 44942 29038 44994
rect 29090 44942 29102 44994
rect 15934 44930 15986 44942
rect 28030 44930 28082 44942
rect 29934 44930 29986 44942
rect 32062 44994 32114 45006
rect 32062 44930 32114 44942
rect 11678 44882 11730 44894
rect 11678 44818 11730 44830
rect 18286 44882 18338 44894
rect 18286 44818 18338 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 14254 44546 14306 44558
rect 14254 44482 14306 44494
rect 3726 44434 3778 44446
rect 3726 44370 3778 44382
rect 4174 44434 4226 44446
rect 20526 44434 20578 44446
rect 25230 44434 25282 44446
rect 9426 44382 9438 44434
rect 9490 44382 9502 44434
rect 9986 44382 9998 44434
rect 10050 44382 10062 44434
rect 12114 44382 12126 44434
rect 12178 44382 12190 44434
rect 15810 44382 15822 44434
rect 15874 44382 15886 44434
rect 19618 44382 19630 44434
rect 19682 44382 19694 44434
rect 24546 44382 24558 44434
rect 24610 44382 24622 44434
rect 4174 44370 4226 44382
rect 20526 44370 20578 44382
rect 25230 44370 25282 44382
rect 30830 44434 30882 44446
rect 30830 44370 30882 44382
rect 31726 44434 31778 44446
rect 31726 44370 31778 44382
rect 32174 44434 32226 44446
rect 32174 44370 32226 44382
rect 15934 44322 15986 44334
rect 20302 44322 20354 44334
rect 26798 44322 26850 44334
rect 3042 44270 3054 44322
rect 3106 44270 3118 44322
rect 6514 44270 6526 44322
rect 6578 44270 6590 44322
rect 12898 44270 12910 44322
rect 12962 44270 12974 44322
rect 15586 44270 15598 44322
rect 15650 44270 15662 44322
rect 16818 44270 16830 44322
rect 16882 44270 16894 44322
rect 21634 44270 21646 44322
rect 21698 44270 21710 44322
rect 15934 44258 15986 44270
rect 20302 44258 20354 44270
rect 26798 44258 26850 44270
rect 27358 44322 27410 44334
rect 29934 44322 29986 44334
rect 28354 44270 28366 44322
rect 28418 44270 28430 44322
rect 27358 44258 27410 44270
rect 29934 44258 29986 44270
rect 5854 44210 5906 44222
rect 13694 44210 13746 44222
rect 2146 44158 2158 44210
rect 2210 44158 2222 44210
rect 7298 44158 7310 44210
rect 7362 44158 7374 44210
rect 5854 44146 5906 44158
rect 13694 44146 13746 44158
rect 14366 44210 14418 44222
rect 20862 44210 20914 44222
rect 26238 44210 26290 44222
rect 17490 44158 17502 44210
rect 17554 44158 17566 44210
rect 22418 44158 22430 44210
rect 22482 44158 22494 44210
rect 14366 44146 14418 44158
rect 20862 44146 20914 44158
rect 26238 44146 26290 44158
rect 26574 44210 26626 44222
rect 26574 44146 26626 44158
rect 27694 44210 27746 44222
rect 27694 44146 27746 44158
rect 29486 44210 29538 44222
rect 29486 44146 29538 44158
rect 30382 44210 30434 44222
rect 30382 44146 30434 44158
rect 4622 44098 4674 44110
rect 4622 44034 4674 44046
rect 5070 44098 5122 44110
rect 5070 44034 5122 44046
rect 5966 44098 6018 44110
rect 5966 44034 6018 44046
rect 13918 44098 13970 44110
rect 13918 44034 13970 44046
rect 14142 44098 14194 44110
rect 14142 44034 14194 44046
rect 16270 44098 16322 44110
rect 16270 44034 16322 44046
rect 20414 44098 20466 44110
rect 20414 44034 20466 44046
rect 20638 44098 20690 44110
rect 20638 44034 20690 44046
rect 25118 44098 25170 44110
rect 25118 44034 25170 44046
rect 25342 44098 25394 44110
rect 25342 44034 25394 44046
rect 25566 44098 25618 44110
rect 25566 44034 25618 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 28590 44098 28642 44110
rect 28590 44034 28642 44046
rect 31278 44098 31330 44110
rect 31278 44034 31330 44046
rect 32622 44098 32674 44110
rect 32622 44034 32674 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 3054 43762 3106 43774
rect 3054 43698 3106 43710
rect 4286 43762 4338 43774
rect 4286 43698 4338 43710
rect 4846 43762 4898 43774
rect 4846 43698 4898 43710
rect 5182 43762 5234 43774
rect 5182 43698 5234 43710
rect 5630 43762 5682 43774
rect 5630 43698 5682 43710
rect 6750 43762 6802 43774
rect 6750 43698 6802 43710
rect 9662 43762 9714 43774
rect 9662 43698 9714 43710
rect 9886 43762 9938 43774
rect 9886 43698 9938 43710
rect 25790 43762 25842 43774
rect 25790 43698 25842 43710
rect 30718 43762 30770 43774
rect 30718 43698 30770 43710
rect 31166 43762 31218 43774
rect 31166 43698 31218 43710
rect 7982 43650 8034 43662
rect 7982 43586 8034 43598
rect 8878 43650 8930 43662
rect 24558 43650 24610 43662
rect 11330 43598 11342 43650
rect 11394 43598 11406 43650
rect 8878 43586 8930 43598
rect 24558 43586 24610 43598
rect 24782 43650 24834 43662
rect 24782 43586 24834 43598
rect 24894 43650 24946 43662
rect 24894 43586 24946 43598
rect 26014 43650 26066 43662
rect 26014 43586 26066 43598
rect 28926 43650 28978 43662
rect 28926 43586 28978 43598
rect 31614 43650 31666 43662
rect 31614 43586 31666 43598
rect 9998 43538 10050 43550
rect 25678 43538 25730 43550
rect 10546 43486 10558 43538
rect 10610 43486 10622 43538
rect 16818 43486 16830 43538
rect 16882 43486 16894 43538
rect 17826 43486 17838 43538
rect 17890 43486 17902 43538
rect 24098 43486 24110 43538
rect 24162 43486 24174 43538
rect 9998 43474 10050 43486
rect 25678 43474 25730 43486
rect 26238 43538 26290 43550
rect 26238 43474 26290 43486
rect 26910 43538 26962 43550
rect 27806 43538 27858 43550
rect 27122 43486 27134 43538
rect 27186 43486 27198 43538
rect 26910 43474 26962 43486
rect 27806 43474 27858 43486
rect 28478 43538 28530 43550
rect 28478 43474 28530 43486
rect 29374 43538 29426 43550
rect 29374 43474 29426 43486
rect 3502 43426 3554 43438
rect 3502 43362 3554 43374
rect 3950 43426 4002 43438
rect 3950 43362 4002 43374
rect 6190 43426 6242 43438
rect 6190 43362 6242 43374
rect 7310 43426 7362 43438
rect 27694 43426 27746 43438
rect 8866 43374 8878 43426
rect 8930 43374 8942 43426
rect 13458 43374 13470 43426
rect 13522 43374 13534 43426
rect 14018 43374 14030 43426
rect 14082 43374 14094 43426
rect 16146 43374 16158 43426
rect 16210 43374 16222 43426
rect 18498 43374 18510 43426
rect 18562 43374 18574 43426
rect 20626 43374 20638 43426
rect 20690 43374 20702 43426
rect 21186 43374 21198 43426
rect 21250 43374 21262 43426
rect 23314 43374 23326 43426
rect 23378 43374 23390 43426
rect 7310 43362 7362 43374
rect 27694 43362 27746 43374
rect 28366 43426 28418 43438
rect 28366 43362 28418 43374
rect 29822 43426 29874 43438
rect 29822 43362 29874 43374
rect 30270 43426 30322 43438
rect 30270 43362 30322 43374
rect 7422 43314 7474 43326
rect 7422 43250 7474 43262
rect 8094 43314 8146 43326
rect 8094 43250 8146 43262
rect 8654 43314 8706 43326
rect 8654 43250 8706 43262
rect 26798 43314 26850 43326
rect 26798 43250 26850 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 8766 42978 8818 42990
rect 8766 42914 8818 42926
rect 9438 42978 9490 42990
rect 9438 42914 9490 42926
rect 13918 42978 13970 42990
rect 13918 42914 13970 42926
rect 27022 42978 27074 42990
rect 27022 42914 27074 42926
rect 4510 42866 4562 42878
rect 4510 42802 4562 42814
rect 5070 42866 5122 42878
rect 5070 42802 5122 42814
rect 5742 42866 5794 42878
rect 5742 42802 5794 42814
rect 6638 42866 6690 42878
rect 6638 42802 6690 42814
rect 9326 42866 9378 42878
rect 14142 42866 14194 42878
rect 9986 42814 9998 42866
rect 10050 42814 10062 42866
rect 9326 42802 9378 42814
rect 14142 42802 14194 42814
rect 14478 42866 14530 42878
rect 20750 42866 20802 42878
rect 27134 42866 27186 42878
rect 16594 42814 16606 42866
rect 16658 42814 16670 42866
rect 21634 42814 21646 42866
rect 21698 42814 21710 42866
rect 14478 42802 14530 42814
rect 20750 42802 20802 42814
rect 27134 42802 27186 42814
rect 27582 42866 27634 42878
rect 27582 42802 27634 42814
rect 28478 42866 28530 42878
rect 28478 42802 28530 42814
rect 29934 42866 29986 42878
rect 29934 42802 29986 42814
rect 30382 42866 30434 42878
rect 30382 42802 30434 42814
rect 7086 42754 7138 42766
rect 14366 42754 14418 42766
rect 12898 42702 12910 42754
rect 12962 42702 12974 42754
rect 7086 42690 7138 42702
rect 14366 42690 14418 42702
rect 15262 42754 15314 42766
rect 20862 42754 20914 42766
rect 15698 42702 15710 42754
rect 15762 42702 15774 42754
rect 16034 42702 16046 42754
rect 16098 42702 16110 42754
rect 19506 42702 19518 42754
rect 19570 42702 19582 42754
rect 20066 42702 20078 42754
rect 20130 42702 20142 42754
rect 24546 42702 24558 42754
rect 24610 42702 24622 42754
rect 15262 42690 15314 42702
rect 20862 42690 20914 42702
rect 7982 42642 8034 42654
rect 7982 42578 8034 42590
rect 8654 42642 8706 42654
rect 20526 42642 20578 42654
rect 25118 42642 25170 42654
rect 12114 42590 12126 42642
rect 12178 42590 12190 42642
rect 18722 42590 18734 42642
rect 18786 42590 18798 42642
rect 23762 42590 23774 42642
rect 23826 42590 23838 42642
rect 8654 42578 8706 42590
rect 20526 42578 20578 42590
rect 25118 42578 25170 42590
rect 25566 42642 25618 42654
rect 25566 42578 25618 42590
rect 26462 42642 26514 42654
rect 26462 42578 26514 42590
rect 1822 42530 1874 42542
rect 1822 42466 1874 42478
rect 6190 42530 6242 42542
rect 6190 42466 6242 42478
rect 7534 42530 7586 42542
rect 7534 42466 7586 42478
rect 8094 42530 8146 42542
rect 8094 42466 8146 42478
rect 14590 42530 14642 42542
rect 14590 42466 14642 42478
rect 15374 42530 15426 42542
rect 15374 42466 15426 42478
rect 15486 42530 15538 42542
rect 15486 42466 15538 42478
rect 20638 42530 20690 42542
rect 20638 42466 20690 42478
rect 25006 42530 25058 42542
rect 25006 42466 25058 42478
rect 25342 42530 25394 42542
rect 25342 42466 25394 42478
rect 26126 42530 26178 42542
rect 26126 42466 26178 42478
rect 28030 42530 28082 42542
rect 28030 42466 28082 42478
rect 29486 42530 29538 42542
rect 29486 42466 29538 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 5630 42194 5682 42206
rect 5630 42130 5682 42142
rect 8990 42194 9042 42206
rect 8990 42130 9042 42142
rect 10894 42194 10946 42206
rect 10894 42130 10946 42142
rect 6190 41970 6242 41982
rect 6190 41906 6242 41918
rect 7870 41970 7922 41982
rect 7870 41906 7922 41918
rect 10222 41970 10274 41982
rect 10222 41906 10274 41918
rect 10334 41970 10386 41982
rect 25790 41970 25842 41982
rect 28926 41970 28978 41982
rect 14466 41918 14478 41970
rect 14530 41918 14542 41970
rect 14914 41918 14926 41970
rect 14978 41918 14990 41970
rect 16370 41918 16382 41970
rect 16434 41918 16446 41970
rect 16706 41918 16718 41970
rect 16770 41918 16782 41970
rect 20514 41918 20526 41970
rect 20578 41918 20590 41970
rect 24098 41918 24110 41970
rect 24162 41918 24174 41970
rect 25890 41918 25902 41970
rect 25954 41967 25966 41970
rect 26114 41967 26126 41970
rect 25954 41921 26126 41967
rect 25954 41918 25966 41921
rect 26114 41918 26126 41921
rect 26178 41918 26190 41970
rect 10334 41906 10386 41918
rect 25790 41906 25842 41918
rect 28926 41906 28978 41918
rect 29374 41970 29426 41982
rect 29374 41906 29426 41918
rect 5294 41858 5346 41870
rect 5294 41794 5346 41806
rect 6638 41858 6690 41870
rect 6638 41794 6690 41806
rect 7086 41858 7138 41870
rect 7086 41794 7138 41806
rect 7422 41858 7474 41870
rect 7422 41794 7474 41806
rect 8318 41858 8370 41870
rect 8318 41794 8370 41806
rect 9662 41858 9714 41870
rect 9662 41794 9714 41806
rect 11454 41858 11506 41870
rect 16942 41858 16994 41870
rect 24782 41858 24834 41870
rect 12002 41806 12014 41858
rect 12066 41806 12078 41858
rect 17714 41806 17726 41858
rect 17778 41806 17790 41858
rect 19842 41806 19854 41858
rect 19906 41806 19918 41858
rect 21186 41806 21198 41858
rect 21250 41806 21262 41858
rect 23314 41806 23326 41858
rect 23378 41806 23390 41858
rect 11454 41794 11506 41806
rect 16942 41794 16994 41806
rect 24782 41794 24834 41806
rect 26238 41858 26290 41870
rect 26238 41794 26290 41806
rect 26686 41858 26738 41870
rect 26686 41794 26738 41806
rect 27134 41858 27186 41870
rect 27134 41794 27186 41806
rect 27582 41858 27634 41870
rect 27582 41794 27634 41806
rect 28030 41858 28082 41870
rect 28030 41794 28082 41806
rect 28478 41858 28530 41870
rect 28478 41794 28530 41806
rect 24670 41746 24722 41758
rect 5282 41694 5294 41746
rect 5346 41743 5358 41746
rect 5842 41743 5854 41746
rect 5346 41697 5854 41743
rect 5346 41694 5358 41697
rect 5842 41694 5854 41697
rect 5906 41743 5918 41746
rect 6738 41743 6750 41746
rect 5906 41697 6750 41743
rect 5906 41694 5918 41697
rect 6738 41694 6750 41697
rect 6802 41694 6814 41746
rect 7858 41694 7870 41746
rect 7922 41743 7934 41746
rect 8306 41743 8318 41746
rect 7922 41697 8318 41743
rect 7922 41694 7934 41697
rect 8306 41694 8318 41697
rect 8370 41694 8382 41746
rect 24670 41682 24722 41694
rect 25678 41746 25730 41758
rect 27010 41694 27022 41746
rect 27074 41743 27086 41746
rect 27570 41743 27582 41746
rect 27074 41697 27582 41743
rect 27074 41694 27086 41697
rect 27570 41694 27582 41697
rect 27634 41694 27646 41746
rect 25678 41682 25730 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 15486 41410 15538 41422
rect 7410 41358 7422 41410
rect 7474 41407 7486 41410
rect 8418 41407 8430 41410
rect 7474 41361 8430 41407
rect 7474 41358 7486 41361
rect 8418 41358 8430 41361
rect 8482 41358 8494 41410
rect 15486 41346 15538 41358
rect 15598 41410 15650 41422
rect 15598 41346 15650 41358
rect 15822 41410 15874 41422
rect 25554 41358 25566 41410
rect 25618 41407 25630 41410
rect 26674 41407 26686 41410
rect 25618 41361 26686 41407
rect 25618 41358 25630 41361
rect 26674 41358 26686 41361
rect 26738 41358 26750 41410
rect 15822 41346 15874 41358
rect 6414 41298 6466 41310
rect 6414 41234 6466 41246
rect 7310 41298 7362 41310
rect 7310 41234 7362 41246
rect 7758 41298 7810 41310
rect 7758 41234 7810 41246
rect 8094 41298 8146 41310
rect 8094 41234 8146 41246
rect 8654 41298 8706 41310
rect 8654 41234 8706 41246
rect 9550 41298 9602 41310
rect 24782 41298 24834 41310
rect 10770 41246 10782 41298
rect 10834 41246 10846 41298
rect 12898 41246 12910 41298
rect 12962 41246 12974 41298
rect 16594 41246 16606 41298
rect 16658 41246 16670 41298
rect 18722 41246 18734 41298
rect 18786 41246 18798 41298
rect 9550 41234 9602 41246
rect 24782 41234 24834 41246
rect 25342 41298 25394 41310
rect 25342 41234 25394 41246
rect 26686 41298 26738 41310
rect 26686 41234 26738 41246
rect 27246 41298 27298 41310
rect 27246 41234 27298 41246
rect 27694 41298 27746 41310
rect 27694 41234 27746 41246
rect 28030 41298 28082 41310
rect 28030 41234 28082 41246
rect 9102 41186 9154 41198
rect 14254 41186 14306 41198
rect 9986 41134 9998 41186
rect 10050 41134 10062 41186
rect 9102 41122 9154 41134
rect 14254 41122 14306 41134
rect 14702 41186 14754 41198
rect 14702 41122 14754 41134
rect 15934 41186 15986 41198
rect 19966 41186 20018 41198
rect 19506 41134 19518 41186
rect 19570 41134 19582 41186
rect 15934 41122 15986 41134
rect 19966 41122 20018 41134
rect 20414 41186 20466 41198
rect 20414 41122 20466 41134
rect 20526 41186 20578 41198
rect 20526 41122 20578 41134
rect 21646 41186 21698 41198
rect 21646 41122 21698 41134
rect 21758 41186 21810 41198
rect 26238 41186 26290 41198
rect 23202 41134 23214 41186
rect 23266 41134 23278 41186
rect 23986 41134 23998 41186
rect 24050 41134 24062 41186
rect 21758 41122 21810 41134
rect 26238 41122 26290 41134
rect 13806 41074 13858 41086
rect 13806 41010 13858 41022
rect 22094 41074 22146 41086
rect 22094 41010 22146 41022
rect 22766 41074 22818 41086
rect 22766 41010 22818 41022
rect 23774 41074 23826 41086
rect 23774 41010 23826 41022
rect 6750 40962 6802 40974
rect 6750 40898 6802 40910
rect 14814 40962 14866 40974
rect 14814 40898 14866 40910
rect 14926 40962 14978 40974
rect 14926 40898 14978 40910
rect 20638 40962 20690 40974
rect 20638 40898 20690 40910
rect 21870 40962 21922 40974
rect 21870 40898 21922 40910
rect 22654 40962 22706 40974
rect 22654 40898 22706 40910
rect 22990 40962 23042 40974
rect 22990 40898 23042 40910
rect 24670 40962 24722 40974
rect 24670 40898 24722 40910
rect 25790 40962 25842 40974
rect 25790 40898 25842 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 7310 40626 7362 40638
rect 7310 40562 7362 40574
rect 7758 40626 7810 40638
rect 7758 40562 7810 40574
rect 8654 40626 8706 40638
rect 8654 40562 8706 40574
rect 9102 40626 9154 40638
rect 9102 40562 9154 40574
rect 10222 40626 10274 40638
rect 10222 40562 10274 40574
rect 10670 40626 10722 40638
rect 10670 40562 10722 40574
rect 11230 40626 11282 40638
rect 11230 40562 11282 40574
rect 15486 40626 15538 40638
rect 15486 40562 15538 40574
rect 16494 40626 16546 40638
rect 16494 40562 16546 40574
rect 21646 40626 21698 40638
rect 21646 40562 21698 40574
rect 22318 40626 22370 40638
rect 22318 40562 22370 40574
rect 23998 40626 24050 40638
rect 23998 40562 24050 40574
rect 24558 40626 24610 40638
rect 24558 40562 24610 40574
rect 25566 40626 25618 40638
rect 25566 40562 25618 40574
rect 26462 40626 26514 40638
rect 26462 40562 26514 40574
rect 26910 40626 26962 40638
rect 26910 40562 26962 40574
rect 27358 40626 27410 40638
rect 27358 40562 27410 40574
rect 11342 40514 11394 40526
rect 11342 40450 11394 40462
rect 15822 40514 15874 40526
rect 15822 40450 15874 40462
rect 16382 40514 16434 40526
rect 16382 40450 16434 40462
rect 16942 40514 16994 40526
rect 21198 40514 21250 40526
rect 19842 40462 19854 40514
rect 19906 40462 19918 40514
rect 16942 40450 16994 40462
rect 21198 40450 21250 40462
rect 22542 40514 22594 40526
rect 22542 40450 22594 40462
rect 24110 40514 24162 40526
rect 24110 40450 24162 40462
rect 48078 40514 48130 40526
rect 48078 40450 48130 40462
rect 8206 40402 8258 40414
rect 16606 40402 16658 40414
rect 21422 40402 21474 40414
rect 14242 40350 14254 40402
rect 14306 40350 14318 40402
rect 14914 40350 14926 40402
rect 14978 40350 14990 40402
rect 20626 40350 20638 40402
rect 20690 40350 20702 40402
rect 8206 40338 8258 40350
rect 16606 40338 16658 40350
rect 21422 40338 21474 40350
rect 21758 40402 21810 40414
rect 21758 40338 21810 40350
rect 22878 40402 22930 40414
rect 22878 40338 22930 40350
rect 26014 40402 26066 40414
rect 26014 40338 26066 40350
rect 9886 40290 9938 40302
rect 23326 40290 23378 40302
rect 11890 40238 11902 40290
rect 11954 40238 11966 40290
rect 17714 40238 17726 40290
rect 17778 40238 17790 40290
rect 9886 40226 9938 40238
rect 23326 40226 23378 40238
rect 22206 40178 22258 40190
rect 6962 40126 6974 40178
rect 7026 40175 7038 40178
rect 8194 40175 8206 40178
rect 7026 40129 8206 40175
rect 7026 40126 7038 40129
rect 8194 40126 8206 40129
rect 8258 40126 8270 40178
rect 8418 40126 8430 40178
rect 8482 40175 8494 40178
rect 9090 40175 9102 40178
rect 8482 40129 9102 40175
rect 8482 40126 8494 40129
rect 9090 40126 9102 40129
rect 9154 40126 9166 40178
rect 22206 40114 22258 40126
rect 23438 40178 23490 40190
rect 23438 40114 23490 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 23090 39790 23102 39842
rect 23154 39839 23166 39842
rect 23314 39839 23326 39842
rect 23154 39793 23326 39839
rect 23154 39790 23166 39793
rect 23314 39790 23326 39793
rect 23378 39790 23390 39842
rect 23538 39790 23550 39842
rect 23602 39839 23614 39842
rect 23874 39839 23886 39842
rect 23602 39793 23886 39839
rect 23602 39790 23614 39793
rect 23874 39790 23886 39793
rect 23938 39839 23950 39842
rect 24434 39839 24446 39842
rect 23938 39793 24446 39839
rect 23938 39790 23950 39793
rect 24434 39790 24446 39793
rect 24498 39790 24510 39842
rect 8318 39730 8370 39742
rect 8318 39666 8370 39678
rect 8766 39730 8818 39742
rect 8766 39666 8818 39678
rect 9102 39730 9154 39742
rect 9102 39666 9154 39678
rect 9550 39730 9602 39742
rect 9550 39666 9602 39678
rect 9998 39730 10050 39742
rect 9998 39666 10050 39678
rect 10558 39730 10610 39742
rect 10558 39666 10610 39678
rect 11454 39730 11506 39742
rect 11454 39666 11506 39678
rect 13694 39730 13746 39742
rect 13694 39666 13746 39678
rect 14254 39730 14306 39742
rect 14254 39666 14306 39678
rect 15710 39730 15762 39742
rect 20302 39730 20354 39742
rect 19282 39678 19294 39730
rect 19346 39678 19358 39730
rect 15710 39666 15762 39678
rect 20302 39666 20354 39678
rect 20862 39730 20914 39742
rect 20862 39666 20914 39678
rect 23550 39730 23602 39742
rect 23550 39666 23602 39678
rect 24446 39730 24498 39742
rect 24446 39666 24498 39678
rect 25006 39730 25058 39742
rect 25006 39666 25058 39678
rect 25342 39730 25394 39742
rect 25342 39666 25394 39678
rect 14142 39618 14194 39630
rect 14142 39554 14194 39566
rect 14814 39618 14866 39630
rect 14814 39554 14866 39566
rect 15598 39618 15650 39630
rect 15598 39554 15650 39566
rect 15822 39618 15874 39630
rect 20190 39618 20242 39630
rect 16370 39566 16382 39618
rect 16434 39566 16446 39618
rect 17154 39566 17166 39618
rect 17218 39566 17230 39618
rect 15822 39554 15874 39566
rect 20190 39554 20242 39566
rect 20414 39618 20466 39630
rect 23998 39618 24050 39630
rect 22754 39566 22766 39618
rect 22818 39615 22830 39618
rect 22978 39615 22990 39618
rect 22818 39569 22990 39615
rect 22818 39566 22830 39569
rect 22978 39566 22990 39569
rect 23042 39566 23054 39618
rect 20414 39554 20466 39566
rect 23998 39554 24050 39566
rect 25790 39618 25842 39630
rect 25790 39554 25842 39566
rect 12014 39506 12066 39518
rect 12014 39442 12066 39454
rect 12910 39506 12962 39518
rect 12910 39442 12962 39454
rect 15262 39506 15314 39518
rect 15262 39442 15314 39454
rect 19966 39506 20018 39518
rect 19966 39442 20018 39454
rect 21646 39506 21698 39518
rect 21646 39442 21698 39454
rect 21982 39506 22034 39518
rect 21982 39442 22034 39454
rect 22542 39506 22594 39518
rect 22542 39442 22594 39454
rect 23102 39506 23154 39518
rect 23102 39442 23154 39454
rect 11006 39394 11058 39406
rect 11006 39330 11058 39342
rect 12574 39394 12626 39406
rect 12574 39330 12626 39342
rect 14366 39394 14418 39406
rect 14366 39330 14418 39342
rect 26238 39394 26290 39406
rect 26238 39330 26290 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 9998 39058 10050 39070
rect 9998 38994 10050 39006
rect 10446 39058 10498 39070
rect 10446 38994 10498 39006
rect 11342 39058 11394 39070
rect 11342 38994 11394 39006
rect 11902 39058 11954 39070
rect 11902 38994 11954 39006
rect 12350 39058 12402 39070
rect 12350 38994 12402 39006
rect 12798 39058 12850 39070
rect 12798 38994 12850 39006
rect 17950 39058 18002 39070
rect 17950 38994 18002 39006
rect 18958 39058 19010 39070
rect 18958 38994 19010 39006
rect 19070 39058 19122 39070
rect 19070 38994 19122 39006
rect 19294 39058 19346 39070
rect 19294 38994 19346 39006
rect 21310 39058 21362 39070
rect 21310 38994 21362 39006
rect 21870 39058 21922 39070
rect 21870 38994 21922 39006
rect 22430 39058 22482 39070
rect 22430 38994 22482 39006
rect 23326 39058 23378 39070
rect 23326 38994 23378 39006
rect 23774 39058 23826 39070
rect 23774 38994 23826 39006
rect 24334 39058 24386 39070
rect 24334 38994 24386 39006
rect 24670 39058 24722 39070
rect 24670 38994 24722 39006
rect 1822 38946 1874 38958
rect 16718 38946 16770 38958
rect 14018 38894 14030 38946
rect 14082 38894 14094 38946
rect 1822 38882 1874 38894
rect 16718 38882 16770 38894
rect 16830 38946 16882 38958
rect 16830 38882 16882 38894
rect 17838 38946 17890 38958
rect 17838 38882 17890 38894
rect 19966 38946 20018 38958
rect 19966 38882 20018 38894
rect 20974 38946 21026 38958
rect 20974 38882 21026 38894
rect 21982 38946 22034 38958
rect 22082 38894 22094 38946
rect 22146 38943 22158 38946
rect 22306 38943 22318 38946
rect 22146 38897 22318 38943
rect 22146 38894 22158 38897
rect 22306 38894 22318 38897
rect 22370 38894 22382 38946
rect 21982 38882 22034 38894
rect 17054 38834 17106 38846
rect 13234 38782 13246 38834
rect 13298 38782 13310 38834
rect 17054 38770 17106 38782
rect 17726 38834 17778 38846
rect 17726 38770 17778 38782
rect 18398 38834 18450 38846
rect 18398 38770 18450 38782
rect 18846 38834 18898 38846
rect 22990 38834 23042 38846
rect 20178 38782 20190 38834
rect 20242 38782 20254 38834
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 18846 38770 18898 38782
rect 22990 38770 23042 38782
rect 10894 38722 10946 38734
rect 19854 38722 19906 38734
rect 16146 38670 16158 38722
rect 16210 38670 16222 38722
rect 10894 38658 10946 38670
rect 19854 38658 19906 38670
rect 10994 38558 11006 38610
rect 11058 38607 11070 38610
rect 11666 38607 11678 38610
rect 11058 38561 11678 38607
rect 11058 38558 11070 38561
rect 11666 38558 11678 38561
rect 11730 38558 11742 38610
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 12562 38222 12574 38274
rect 12626 38271 12638 38274
rect 13122 38271 13134 38274
rect 12626 38225 13134 38271
rect 12626 38222 12638 38225
rect 13122 38222 13134 38225
rect 13186 38222 13198 38274
rect 20626 38222 20638 38274
rect 20690 38271 20702 38274
rect 21074 38271 21086 38274
rect 20690 38225 21086 38271
rect 20690 38222 20702 38225
rect 21074 38222 21086 38225
rect 21138 38222 21150 38274
rect 10558 38162 10610 38174
rect 10558 38098 10610 38110
rect 11006 38162 11058 38174
rect 11006 38098 11058 38110
rect 12014 38162 12066 38174
rect 12014 38098 12066 38110
rect 12574 38162 12626 38174
rect 12574 38098 12626 38110
rect 13022 38162 13074 38174
rect 13022 38098 13074 38110
rect 14254 38162 14306 38174
rect 21534 38162 21586 38174
rect 18386 38110 18398 38162
rect 18450 38110 18462 38162
rect 14254 38098 14306 38110
rect 21534 38098 21586 38110
rect 22094 38162 22146 38174
rect 22094 38098 22146 38110
rect 22430 38162 22482 38174
rect 22430 38098 22482 38110
rect 22990 38162 23042 38174
rect 22990 38098 23042 38110
rect 24334 38162 24386 38174
rect 24334 38098 24386 38110
rect 18958 38050 19010 38062
rect 15474 37998 15486 38050
rect 15538 37998 15550 38050
rect 18958 37986 19010 37998
rect 20078 38050 20130 38062
rect 20078 37986 20130 37998
rect 23438 38050 23490 38062
rect 23438 37986 23490 37998
rect 14814 37938 14866 37950
rect 14814 37874 14866 37886
rect 14926 37938 14978 37950
rect 19406 37938 19458 37950
rect 16258 37886 16270 37938
rect 16322 37886 16334 37938
rect 14926 37874 14978 37886
rect 19406 37874 19458 37886
rect 20414 37938 20466 37950
rect 20414 37874 20466 37886
rect 13918 37826 13970 37838
rect 13918 37762 13970 37774
rect 19070 37826 19122 37838
rect 19070 37762 19122 37774
rect 19182 37826 19234 37838
rect 19182 37762 19234 37774
rect 20862 37826 20914 37838
rect 20862 37762 20914 37774
rect 23774 37826 23826 37838
rect 23774 37762 23826 37774
rect 48078 37826 48130 37838
rect 48078 37762 48130 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 13134 37490 13186 37502
rect 13134 37426 13186 37438
rect 14142 37490 14194 37502
rect 14142 37426 14194 37438
rect 14590 37490 14642 37502
rect 14590 37426 14642 37438
rect 18174 37490 18226 37502
rect 18174 37426 18226 37438
rect 18846 37490 18898 37502
rect 18846 37426 18898 37438
rect 19854 37490 19906 37502
rect 19854 37426 19906 37438
rect 21198 37490 21250 37502
rect 21198 37426 21250 37438
rect 21758 37490 21810 37502
rect 21758 37426 21810 37438
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 22542 37490 22594 37502
rect 22542 37426 22594 37438
rect 22990 37490 23042 37502
rect 22990 37426 23042 37438
rect 1822 37378 1874 37390
rect 1822 37314 1874 37326
rect 16942 37378 16994 37390
rect 16942 37314 16994 37326
rect 18286 37378 18338 37390
rect 18286 37314 18338 37326
rect 19182 37378 19234 37390
rect 19182 37314 19234 37326
rect 15486 37266 15538 37278
rect 15486 37202 15538 37214
rect 16606 37266 16658 37278
rect 16606 37202 16658 37214
rect 17614 37266 17666 37278
rect 17614 37202 17666 37214
rect 18062 37266 18114 37278
rect 18062 37202 18114 37214
rect 13694 37154 13746 37166
rect 13694 37090 13746 37102
rect 14926 37154 14978 37166
rect 14926 37090 14978 37102
rect 15934 37154 15986 37166
rect 15934 37090 15986 37102
rect 19742 37154 19794 37166
rect 19742 37090 19794 37102
rect 20302 37154 20354 37166
rect 20302 37090 20354 37102
rect 20862 37154 20914 37166
rect 20862 37090 20914 37102
rect 16046 37042 16098 37054
rect 14242 36990 14254 37042
rect 14306 37039 14318 37042
rect 14690 37039 14702 37042
rect 14306 36993 14702 37039
rect 14306 36990 14318 36993
rect 14690 36990 14702 36993
rect 14754 36990 14766 37042
rect 16046 36978 16098 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 16606 36706 16658 36718
rect 16606 36642 16658 36654
rect 14702 36594 14754 36606
rect 14702 36530 14754 36542
rect 15598 36594 15650 36606
rect 15598 36530 15650 36542
rect 16158 36594 16210 36606
rect 16158 36530 16210 36542
rect 17502 36594 17554 36606
rect 17502 36530 17554 36542
rect 18958 36594 19010 36606
rect 18958 36530 19010 36542
rect 19406 36594 19458 36606
rect 19406 36530 19458 36542
rect 20414 36594 20466 36606
rect 20414 36530 20466 36542
rect 20974 36594 21026 36606
rect 20974 36530 21026 36542
rect 21534 36594 21586 36606
rect 21534 36530 21586 36542
rect 22094 36594 22146 36606
rect 22094 36530 22146 36542
rect 16718 36482 16770 36494
rect 18510 36482 18562 36494
rect 17266 36430 17278 36482
rect 17330 36430 17342 36482
rect 16718 36418 16770 36430
rect 18510 36418 18562 36430
rect 17614 36370 17666 36382
rect 17614 36306 17666 36318
rect 15150 36258 15202 36270
rect 15150 36194 15202 36206
rect 18174 36258 18226 36270
rect 18174 36194 18226 36206
rect 19966 36258 20018 36270
rect 19966 36194 20018 36206
rect 48078 36258 48130 36270
rect 48078 36194 48130 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 16158 35922 16210 35934
rect 16158 35858 16210 35870
rect 16606 35922 16658 35934
rect 16606 35858 16658 35870
rect 17726 35922 17778 35934
rect 17726 35858 17778 35870
rect 18174 35922 18226 35934
rect 18174 35858 18226 35870
rect 18622 35922 18674 35934
rect 18622 35858 18674 35870
rect 19070 35922 19122 35934
rect 19070 35858 19122 35870
rect 19518 35922 19570 35934
rect 19518 35858 19570 35870
rect 19966 35922 20018 35934
rect 19966 35858 20018 35870
rect 20862 35922 20914 35934
rect 20862 35858 20914 35870
rect 1822 35810 1874 35822
rect 1822 35746 1874 35758
rect 17054 35698 17106 35710
rect 17054 35634 17106 35646
rect 20414 35586 20466 35598
rect 20414 35522 20466 35534
rect 19506 35422 19518 35474
rect 19570 35471 19582 35474
rect 20402 35471 20414 35474
rect 19570 35425 20414 35471
rect 19570 35422 19582 35425
rect 20402 35422 20414 35425
rect 20466 35422 20478 35474
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 17502 35026 17554 35038
rect 17502 34962 17554 34974
rect 17950 35026 18002 35038
rect 17950 34962 18002 34974
rect 18622 35026 18674 35038
rect 18622 34962 18674 34974
rect 19070 35026 19122 35038
rect 19070 34962 19122 34974
rect 48078 34690 48130 34702
rect 48078 34626 48130 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 1822 33122 1874 33134
rect 1822 33058 1874 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 48078 32674 48130 32686
rect 48078 32610 48130 32622
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 48078 31554 48130 31566
rect 48078 31490 48130 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 1822 29986 1874 29998
rect 1822 29922 1874 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 48078 29538 48130 29550
rect 48078 29474 48130 29486
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 1822 28418 1874 28430
rect 1822 28354 1874 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 1822 26850 1874 26862
rect 1822 26786 1874 26798
rect 48078 26850 48130 26862
rect 48078 26786 48130 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 1822 24834 1874 24846
rect 1822 24770 1874 24782
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 48078 23714 48130 23726
rect 48078 23650 48130 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 3502 23378 3554 23390
rect 3502 23314 3554 23326
rect 3042 23102 3054 23154
rect 3106 23102 3118 23154
rect 2034 22990 2046 23042
rect 2098 22990 2110 23042
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 48078 22146 48130 22158
rect 48078 22082 48130 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 1822 21698 1874 21710
rect 1822 21634 1874 21646
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 1822 19010 1874 19022
rect 1822 18946 1874 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 48078 18562 48130 18574
rect 48078 18498 48130 18510
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 1822 17554 1874 17566
rect 1822 17490 1874 17502
rect 48078 17442 48130 17454
rect 48078 17378 48130 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 1822 15874 1874 15886
rect 1822 15810 1874 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 1822 14306 1874 14318
rect 1822 14242 1874 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 48078 12850 48130 12862
rect 48078 12786 48130 12798
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 48078 12290 48130 12302
rect 48078 12226 48130 12238
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 1822 10722 1874 10734
rect 1822 10658 1874 10670
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 48078 9602 48130 9614
rect 48078 9538 48130 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 1822 9154 1874 9166
rect 1822 9090 1874 9102
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 48078 8034 48130 8046
rect 48078 7970 48130 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 1822 7586 1874 7598
rect 1822 7522 1874 7534
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 48078 6466 48130 6478
rect 48078 6402 48130 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 1822 4450 1874 4462
rect 1822 4386 1874 4398
rect 2494 4450 2546 4462
rect 2494 4386 2546 4398
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 4286 3666 4338 3678
rect 4286 3602 4338 3614
rect 2146 3502 2158 3554
rect 2210 3502 2222 3554
rect 3042 3502 3054 3554
rect 3106 3502 3118 3554
rect 3614 3330 3666 3342
rect 3614 3266 3666 3278
rect 5742 3330 5794 3342
rect 5742 3266 5794 3278
rect 9662 3330 9714 3342
rect 9662 3266 9714 3278
rect 14366 3330 14418 3342
rect 14366 3266 14418 3278
rect 15710 3330 15762 3342
rect 15710 3266 15762 3278
rect 17726 3330 17778 3342
rect 17726 3266 17778 3278
rect 21422 3330 21474 3342
rect 21422 3266 21474 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 29262 3330 29314 3342
rect 29262 3266 29314 3278
rect 31838 3330 31890 3342
rect 31838 3266 31890 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 38558 3330 38610 3342
rect 38558 3266 38610 3278
rect 41022 3330 41074 3342
rect 41022 3266 41074 3278
rect 42590 3330 42642 3342
rect 42590 3266 42642 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 45950 3330 46002 3342
rect 45950 3266 46002 3278
rect 47406 3330 47458 3342
rect 47406 3266 47458 3278
rect 48078 3330 48130 3342
rect 48078 3266 48130 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
rect 40338 1822 40350 1874
rect 40402 1871 40414 1874
rect 41010 1871 41022 1874
rect 40402 1825 41022 1871
rect 40402 1822 40414 1825
rect 41010 1822 41022 1825
rect 41074 1822 41086 1874
rect 8754 1710 8766 1762
rect 8818 1759 8830 1762
rect 9650 1759 9662 1762
rect 8818 1713 9662 1759
rect 8818 1710 8830 1713
rect 9650 1710 9662 1713
rect 9714 1710 9726 1762
rect 20850 1710 20862 1762
rect 20914 1759 20926 1762
rect 21410 1759 21422 1762
rect 20914 1713 21422 1759
rect 20914 1710 20926 1713
rect 21410 1710 21422 1713
rect 21474 1710 21486 1762
<< via1 >>
rect 11902 47854 11954 47906
rect 12798 47854 12850 47906
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 4062 45950 4114 46002
rect 5966 45950 6018 46002
rect 12798 45950 12850 46002
rect 24446 45950 24498 46002
rect 25342 45950 25394 46002
rect 27470 45950 27522 46002
rect 32398 45950 32450 46002
rect 33854 45950 33906 46002
rect 35758 45950 35810 46002
rect 42478 45950 42530 46002
rect 43710 45950 43762 46002
rect 4958 45838 5010 45890
rect 8766 45838 8818 45890
rect 9998 45838 10050 45890
rect 13582 45838 13634 45890
rect 15934 45838 15986 45890
rect 16494 45838 16546 45890
rect 19966 45838 20018 45890
rect 20638 45838 20690 45890
rect 21310 45838 21362 45890
rect 22094 45838 22146 45890
rect 28254 45838 28306 45890
rect 31390 45838 31442 45890
rect 31950 45838 32002 45890
rect 33182 45838 33234 45890
rect 35086 45838 35138 45890
rect 42926 45838 42978 45890
rect 2270 45726 2322 45778
rect 2942 45726 2994 45778
rect 8094 45726 8146 45778
rect 10670 45726 10722 45778
rect 29262 45726 29314 45778
rect 29486 45726 29538 45778
rect 29822 45726 29874 45778
rect 30382 45726 30434 45778
rect 31166 45726 31218 45778
rect 37886 45726 37938 45778
rect 39902 45726 39954 45778
rect 48078 45726 48130 45778
rect 1822 45614 1874 45666
rect 17502 45614 17554 45666
rect 29598 45614 29650 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 1822 45278 1874 45330
rect 2494 45278 2546 45330
rect 3166 45278 3218 45330
rect 3502 45278 3554 45330
rect 5518 45278 5570 45330
rect 12238 45278 12290 45330
rect 23774 45278 23826 45330
rect 24446 45278 24498 45330
rect 26238 45278 26290 45330
rect 27022 45278 27074 45330
rect 30718 45278 30770 45330
rect 31166 45278 31218 45330
rect 33518 45278 33570 45330
rect 34750 45278 34802 45330
rect 6862 45166 6914 45218
rect 18398 45166 18450 45218
rect 27134 45166 27186 45218
rect 27358 45166 27410 45218
rect 29150 45166 29202 45218
rect 29374 45166 29426 45218
rect 30046 45166 30098 45218
rect 30606 45166 30658 45218
rect 31614 45166 31666 45218
rect 6190 45054 6242 45106
rect 9774 45054 9826 45106
rect 10110 45054 10162 45106
rect 10334 45054 10386 45106
rect 11006 45054 11058 45106
rect 11118 45054 11170 45106
rect 11230 45054 11282 45106
rect 14590 45054 14642 45106
rect 15374 45054 15426 45106
rect 16382 45054 16434 45106
rect 17726 45054 17778 45106
rect 17950 45054 18002 45106
rect 18174 45054 18226 45106
rect 18958 45054 19010 45106
rect 20862 45054 20914 45106
rect 21422 45054 21474 45106
rect 24222 45054 24274 45106
rect 24558 45054 24610 45106
rect 24782 45054 24834 45106
rect 25566 45054 25618 45106
rect 26014 45054 26066 45106
rect 26126 45054 26178 45106
rect 26686 45054 26738 45106
rect 27918 45054 27970 45106
rect 28142 45054 28194 45106
rect 28478 45054 28530 45106
rect 32510 45054 32562 45106
rect 4062 44942 4114 44994
rect 4510 44942 4562 44994
rect 4958 44942 5010 44994
rect 5406 44942 5458 44994
rect 8990 44942 9042 44994
rect 10222 44942 10274 44994
rect 11454 44942 11506 44994
rect 15934 44942 15986 44994
rect 16270 44942 16322 44994
rect 19966 44942 20018 44994
rect 28030 44942 28082 44994
rect 29038 44942 29090 44994
rect 29934 44942 29986 44994
rect 32062 44942 32114 44994
rect 11678 44830 11730 44882
rect 18286 44830 18338 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 14254 44494 14306 44546
rect 3726 44382 3778 44434
rect 4174 44382 4226 44434
rect 9438 44382 9490 44434
rect 9998 44382 10050 44434
rect 12126 44382 12178 44434
rect 15822 44382 15874 44434
rect 19630 44382 19682 44434
rect 20526 44382 20578 44434
rect 24558 44382 24610 44434
rect 25230 44382 25282 44434
rect 30830 44382 30882 44434
rect 31726 44382 31778 44434
rect 32174 44382 32226 44434
rect 3054 44270 3106 44322
rect 6526 44270 6578 44322
rect 12910 44270 12962 44322
rect 15598 44270 15650 44322
rect 15934 44270 15986 44322
rect 16830 44270 16882 44322
rect 20302 44270 20354 44322
rect 21646 44270 21698 44322
rect 26798 44270 26850 44322
rect 27358 44270 27410 44322
rect 28366 44270 28418 44322
rect 29934 44270 29986 44322
rect 2158 44158 2210 44210
rect 5854 44158 5906 44210
rect 7310 44158 7362 44210
rect 13694 44158 13746 44210
rect 14366 44158 14418 44210
rect 17502 44158 17554 44210
rect 20862 44158 20914 44210
rect 22430 44158 22482 44210
rect 26238 44158 26290 44210
rect 26574 44158 26626 44210
rect 27694 44158 27746 44210
rect 29486 44158 29538 44210
rect 30382 44158 30434 44210
rect 4622 44046 4674 44098
rect 5070 44046 5122 44098
rect 5966 44046 6018 44098
rect 13918 44046 13970 44098
rect 14142 44046 14194 44098
rect 16270 44046 16322 44098
rect 20414 44046 20466 44098
rect 20638 44046 20690 44098
rect 25118 44046 25170 44098
rect 25342 44046 25394 44098
rect 25566 44046 25618 44098
rect 26462 44046 26514 44098
rect 28590 44046 28642 44098
rect 31278 44046 31330 44098
rect 32622 44046 32674 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 3054 43710 3106 43762
rect 4286 43710 4338 43762
rect 4846 43710 4898 43762
rect 5182 43710 5234 43762
rect 5630 43710 5682 43762
rect 6750 43710 6802 43762
rect 9662 43710 9714 43762
rect 9886 43710 9938 43762
rect 25790 43710 25842 43762
rect 30718 43710 30770 43762
rect 31166 43710 31218 43762
rect 7982 43598 8034 43650
rect 8878 43598 8930 43650
rect 11342 43598 11394 43650
rect 24558 43598 24610 43650
rect 24782 43598 24834 43650
rect 24894 43598 24946 43650
rect 26014 43598 26066 43650
rect 28926 43598 28978 43650
rect 31614 43598 31666 43650
rect 9998 43486 10050 43538
rect 10558 43486 10610 43538
rect 16830 43486 16882 43538
rect 17838 43486 17890 43538
rect 24110 43486 24162 43538
rect 25678 43486 25730 43538
rect 26238 43486 26290 43538
rect 26910 43486 26962 43538
rect 27134 43486 27186 43538
rect 27806 43486 27858 43538
rect 28478 43486 28530 43538
rect 29374 43486 29426 43538
rect 3502 43374 3554 43426
rect 3950 43374 4002 43426
rect 6190 43374 6242 43426
rect 7310 43374 7362 43426
rect 8878 43374 8930 43426
rect 13470 43374 13522 43426
rect 14030 43374 14082 43426
rect 16158 43374 16210 43426
rect 18510 43374 18562 43426
rect 20638 43374 20690 43426
rect 21198 43374 21250 43426
rect 23326 43374 23378 43426
rect 27694 43374 27746 43426
rect 28366 43374 28418 43426
rect 29822 43374 29874 43426
rect 30270 43374 30322 43426
rect 7422 43262 7474 43314
rect 8094 43262 8146 43314
rect 8654 43262 8706 43314
rect 26798 43262 26850 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 8766 42926 8818 42978
rect 9438 42926 9490 42978
rect 13918 42926 13970 42978
rect 27022 42926 27074 42978
rect 4510 42814 4562 42866
rect 5070 42814 5122 42866
rect 5742 42814 5794 42866
rect 6638 42814 6690 42866
rect 9326 42814 9378 42866
rect 9998 42814 10050 42866
rect 14142 42814 14194 42866
rect 14478 42814 14530 42866
rect 16606 42814 16658 42866
rect 20750 42814 20802 42866
rect 21646 42814 21698 42866
rect 27134 42814 27186 42866
rect 27582 42814 27634 42866
rect 28478 42814 28530 42866
rect 29934 42814 29986 42866
rect 30382 42814 30434 42866
rect 7086 42702 7138 42754
rect 12910 42702 12962 42754
rect 14366 42702 14418 42754
rect 15262 42702 15314 42754
rect 15710 42702 15762 42754
rect 16046 42702 16098 42754
rect 19518 42702 19570 42754
rect 20078 42702 20130 42754
rect 20862 42702 20914 42754
rect 24558 42702 24610 42754
rect 7982 42590 8034 42642
rect 8654 42590 8706 42642
rect 12126 42590 12178 42642
rect 18734 42590 18786 42642
rect 20526 42590 20578 42642
rect 23774 42590 23826 42642
rect 25118 42590 25170 42642
rect 25566 42590 25618 42642
rect 26462 42590 26514 42642
rect 1822 42478 1874 42530
rect 6190 42478 6242 42530
rect 7534 42478 7586 42530
rect 8094 42478 8146 42530
rect 14590 42478 14642 42530
rect 15374 42478 15426 42530
rect 15486 42478 15538 42530
rect 20638 42478 20690 42530
rect 25006 42478 25058 42530
rect 25342 42478 25394 42530
rect 26126 42478 26178 42530
rect 28030 42478 28082 42530
rect 29486 42478 29538 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 5630 42142 5682 42194
rect 8990 42142 9042 42194
rect 10894 42142 10946 42194
rect 6190 41918 6242 41970
rect 7870 41918 7922 41970
rect 10222 41918 10274 41970
rect 10334 41918 10386 41970
rect 14478 41918 14530 41970
rect 14926 41918 14978 41970
rect 16382 41918 16434 41970
rect 16718 41918 16770 41970
rect 20526 41918 20578 41970
rect 24110 41918 24162 41970
rect 25790 41918 25842 41970
rect 25902 41918 25954 41970
rect 26126 41918 26178 41970
rect 28926 41918 28978 41970
rect 29374 41918 29426 41970
rect 5294 41806 5346 41858
rect 6638 41806 6690 41858
rect 7086 41806 7138 41858
rect 7422 41806 7474 41858
rect 8318 41806 8370 41858
rect 9662 41806 9714 41858
rect 11454 41806 11506 41858
rect 12014 41806 12066 41858
rect 16942 41806 16994 41858
rect 17726 41806 17778 41858
rect 19854 41806 19906 41858
rect 21198 41806 21250 41858
rect 23326 41806 23378 41858
rect 24782 41806 24834 41858
rect 26238 41806 26290 41858
rect 26686 41806 26738 41858
rect 27134 41806 27186 41858
rect 27582 41806 27634 41858
rect 28030 41806 28082 41858
rect 28478 41806 28530 41858
rect 5294 41694 5346 41746
rect 5854 41694 5906 41746
rect 6750 41694 6802 41746
rect 7870 41694 7922 41746
rect 8318 41694 8370 41746
rect 24670 41694 24722 41746
rect 25678 41694 25730 41746
rect 27022 41694 27074 41746
rect 27582 41694 27634 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 7422 41358 7474 41410
rect 8430 41358 8482 41410
rect 15486 41358 15538 41410
rect 15598 41358 15650 41410
rect 15822 41358 15874 41410
rect 25566 41358 25618 41410
rect 26686 41358 26738 41410
rect 6414 41246 6466 41298
rect 7310 41246 7362 41298
rect 7758 41246 7810 41298
rect 8094 41246 8146 41298
rect 8654 41246 8706 41298
rect 9550 41246 9602 41298
rect 10782 41246 10834 41298
rect 12910 41246 12962 41298
rect 16606 41246 16658 41298
rect 18734 41246 18786 41298
rect 24782 41246 24834 41298
rect 25342 41246 25394 41298
rect 26686 41246 26738 41298
rect 27246 41246 27298 41298
rect 27694 41246 27746 41298
rect 28030 41246 28082 41298
rect 9102 41134 9154 41186
rect 9998 41134 10050 41186
rect 14254 41134 14306 41186
rect 14702 41134 14754 41186
rect 15934 41134 15986 41186
rect 19518 41134 19570 41186
rect 19966 41134 20018 41186
rect 20414 41134 20466 41186
rect 20526 41134 20578 41186
rect 21646 41134 21698 41186
rect 21758 41134 21810 41186
rect 23214 41134 23266 41186
rect 23998 41134 24050 41186
rect 26238 41134 26290 41186
rect 13806 41022 13858 41074
rect 22094 41022 22146 41074
rect 22766 41022 22818 41074
rect 23774 41022 23826 41074
rect 6750 40910 6802 40962
rect 14814 40910 14866 40962
rect 14926 40910 14978 40962
rect 20638 40910 20690 40962
rect 21870 40910 21922 40962
rect 22654 40910 22706 40962
rect 22990 40910 23042 40962
rect 24670 40910 24722 40962
rect 25790 40910 25842 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 7310 40574 7362 40626
rect 7758 40574 7810 40626
rect 8654 40574 8706 40626
rect 9102 40574 9154 40626
rect 10222 40574 10274 40626
rect 10670 40574 10722 40626
rect 11230 40574 11282 40626
rect 15486 40574 15538 40626
rect 16494 40574 16546 40626
rect 21646 40574 21698 40626
rect 22318 40574 22370 40626
rect 23998 40574 24050 40626
rect 24558 40574 24610 40626
rect 25566 40574 25618 40626
rect 26462 40574 26514 40626
rect 26910 40574 26962 40626
rect 27358 40574 27410 40626
rect 11342 40462 11394 40514
rect 15822 40462 15874 40514
rect 16382 40462 16434 40514
rect 16942 40462 16994 40514
rect 19854 40462 19906 40514
rect 21198 40462 21250 40514
rect 22542 40462 22594 40514
rect 24110 40462 24162 40514
rect 48078 40462 48130 40514
rect 8206 40350 8258 40402
rect 14254 40350 14306 40402
rect 14926 40350 14978 40402
rect 16606 40350 16658 40402
rect 20638 40350 20690 40402
rect 21422 40350 21474 40402
rect 21758 40350 21810 40402
rect 22878 40350 22930 40402
rect 26014 40350 26066 40402
rect 9886 40238 9938 40290
rect 11902 40238 11954 40290
rect 17726 40238 17778 40290
rect 23326 40238 23378 40290
rect 6974 40126 7026 40178
rect 8206 40126 8258 40178
rect 8430 40126 8482 40178
rect 9102 40126 9154 40178
rect 22206 40126 22258 40178
rect 23438 40126 23490 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 23102 39790 23154 39842
rect 23326 39790 23378 39842
rect 23550 39790 23602 39842
rect 23886 39790 23938 39842
rect 24446 39790 24498 39842
rect 8318 39678 8370 39730
rect 8766 39678 8818 39730
rect 9102 39678 9154 39730
rect 9550 39678 9602 39730
rect 9998 39678 10050 39730
rect 10558 39678 10610 39730
rect 11454 39678 11506 39730
rect 13694 39678 13746 39730
rect 14254 39678 14306 39730
rect 15710 39678 15762 39730
rect 19294 39678 19346 39730
rect 20302 39678 20354 39730
rect 20862 39678 20914 39730
rect 23550 39678 23602 39730
rect 24446 39678 24498 39730
rect 25006 39678 25058 39730
rect 25342 39678 25394 39730
rect 14142 39566 14194 39618
rect 14814 39566 14866 39618
rect 15598 39566 15650 39618
rect 15822 39566 15874 39618
rect 16382 39566 16434 39618
rect 17166 39566 17218 39618
rect 20190 39566 20242 39618
rect 20414 39566 20466 39618
rect 22766 39566 22818 39618
rect 22990 39566 23042 39618
rect 23998 39566 24050 39618
rect 25790 39566 25842 39618
rect 12014 39454 12066 39506
rect 12910 39454 12962 39506
rect 15262 39454 15314 39506
rect 19966 39454 20018 39506
rect 21646 39454 21698 39506
rect 21982 39454 22034 39506
rect 22542 39454 22594 39506
rect 23102 39454 23154 39506
rect 11006 39342 11058 39394
rect 12574 39342 12626 39394
rect 14366 39342 14418 39394
rect 26238 39342 26290 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 9998 39006 10050 39058
rect 10446 39006 10498 39058
rect 11342 39006 11394 39058
rect 11902 39006 11954 39058
rect 12350 39006 12402 39058
rect 12798 39006 12850 39058
rect 17950 39006 18002 39058
rect 18958 39006 19010 39058
rect 19070 39006 19122 39058
rect 19294 39006 19346 39058
rect 21310 39006 21362 39058
rect 21870 39006 21922 39058
rect 22430 39006 22482 39058
rect 23326 39006 23378 39058
rect 23774 39006 23826 39058
rect 24334 39006 24386 39058
rect 24670 39006 24722 39058
rect 1822 38894 1874 38946
rect 14030 38894 14082 38946
rect 16718 38894 16770 38946
rect 16830 38894 16882 38946
rect 17838 38894 17890 38946
rect 19966 38894 20018 38946
rect 20974 38894 21026 38946
rect 21982 38894 22034 38946
rect 22094 38894 22146 38946
rect 22318 38894 22370 38946
rect 13246 38782 13298 38834
rect 17054 38782 17106 38834
rect 17726 38782 17778 38834
rect 18398 38782 18450 38834
rect 18846 38782 18898 38834
rect 20190 38782 20242 38834
rect 20414 38782 20466 38834
rect 22990 38782 23042 38834
rect 10894 38670 10946 38722
rect 16158 38670 16210 38722
rect 19854 38670 19906 38722
rect 11006 38558 11058 38610
rect 11678 38558 11730 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 12574 38222 12626 38274
rect 13134 38222 13186 38274
rect 20638 38222 20690 38274
rect 21086 38222 21138 38274
rect 10558 38110 10610 38162
rect 11006 38110 11058 38162
rect 12014 38110 12066 38162
rect 12574 38110 12626 38162
rect 13022 38110 13074 38162
rect 14254 38110 14306 38162
rect 18398 38110 18450 38162
rect 21534 38110 21586 38162
rect 22094 38110 22146 38162
rect 22430 38110 22482 38162
rect 22990 38110 23042 38162
rect 24334 38110 24386 38162
rect 15486 37998 15538 38050
rect 18958 37998 19010 38050
rect 20078 37998 20130 38050
rect 23438 37998 23490 38050
rect 14814 37886 14866 37938
rect 14926 37886 14978 37938
rect 16270 37886 16322 37938
rect 19406 37886 19458 37938
rect 20414 37886 20466 37938
rect 13918 37774 13970 37826
rect 19070 37774 19122 37826
rect 19182 37774 19234 37826
rect 20862 37774 20914 37826
rect 23774 37774 23826 37826
rect 48078 37774 48130 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 13134 37438 13186 37490
rect 14142 37438 14194 37490
rect 14590 37438 14642 37490
rect 18174 37438 18226 37490
rect 18846 37438 18898 37490
rect 19854 37438 19906 37490
rect 21198 37438 21250 37490
rect 21758 37438 21810 37490
rect 22094 37438 22146 37490
rect 22542 37438 22594 37490
rect 22990 37438 23042 37490
rect 1822 37326 1874 37378
rect 16942 37326 16994 37378
rect 18286 37326 18338 37378
rect 19182 37326 19234 37378
rect 15486 37214 15538 37266
rect 16606 37214 16658 37266
rect 17614 37214 17666 37266
rect 18062 37214 18114 37266
rect 13694 37102 13746 37154
rect 14926 37102 14978 37154
rect 15934 37102 15986 37154
rect 19742 37102 19794 37154
rect 20302 37102 20354 37154
rect 20862 37102 20914 37154
rect 14254 36990 14306 37042
rect 14702 36990 14754 37042
rect 16046 36990 16098 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 16606 36654 16658 36706
rect 14702 36542 14754 36594
rect 15598 36542 15650 36594
rect 16158 36542 16210 36594
rect 17502 36542 17554 36594
rect 18958 36542 19010 36594
rect 19406 36542 19458 36594
rect 20414 36542 20466 36594
rect 20974 36542 21026 36594
rect 21534 36542 21586 36594
rect 22094 36542 22146 36594
rect 16718 36430 16770 36482
rect 17278 36430 17330 36482
rect 18510 36430 18562 36482
rect 17614 36318 17666 36370
rect 15150 36206 15202 36258
rect 18174 36206 18226 36258
rect 19966 36206 20018 36258
rect 48078 36206 48130 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 16158 35870 16210 35922
rect 16606 35870 16658 35922
rect 17726 35870 17778 35922
rect 18174 35870 18226 35922
rect 18622 35870 18674 35922
rect 19070 35870 19122 35922
rect 19518 35870 19570 35922
rect 19966 35870 20018 35922
rect 20862 35870 20914 35922
rect 1822 35758 1874 35810
rect 17054 35646 17106 35698
rect 20414 35534 20466 35586
rect 19518 35422 19570 35474
rect 20414 35422 20466 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 17502 34974 17554 35026
rect 17950 34974 18002 35026
rect 18622 34974 18674 35026
rect 19070 34974 19122 35026
rect 48078 34638 48130 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 1822 33070 1874 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 48078 32622 48130 32674
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 48078 31502 48130 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 1822 29934 1874 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 48078 29486 48130 29538
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 1822 28366 1874 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1822 26798 1874 26850
rect 48078 26798 48130 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 1822 24782 1874 24834
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 48078 23662 48130 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 3502 23326 3554 23378
rect 3054 23102 3106 23154
rect 2046 22990 2098 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 48078 22094 48130 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 1822 21646 1874 21698
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 1822 18958 1874 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 48078 18510 48130 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 1822 17502 1874 17554
rect 48078 17390 48130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 1822 15822 1874 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 1822 14254 1874 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 48078 12798 48130 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 48078 12238 48130 12290
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 1822 10670 1874 10722
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 48078 9550 48130 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 1822 9102 1874 9154
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 48078 7982 48130 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 1822 7534 1874 7586
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 48078 6414 48130 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 1822 4398 1874 4450
rect 2494 4398 2546 4450
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 4286 3614 4338 3666
rect 2158 3502 2210 3554
rect 3054 3502 3106 3554
rect 3614 3278 3666 3330
rect 5742 3278 5794 3330
rect 9662 3278 9714 3330
rect 14366 3278 14418 3330
rect 15710 3278 15762 3330
rect 17726 3278 17778 3330
rect 21422 3278 21474 3330
rect 23102 3278 23154 3330
rect 26462 3278 26514 3330
rect 29262 3278 29314 3330
rect 31838 3278 31890 3330
rect 35198 3278 35250 3330
rect 38558 3278 38610 3330
rect 41022 3278 41074 3330
rect 42590 3278 42642 3330
rect 43934 3278 43986 3330
rect 45950 3278 46002 3330
rect 47406 3278 47458 3330
rect 48078 3278 48130 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 40350 1822 40402 1874
rect 41022 1822 41074 1874
rect 8766 1710 8818 1762
rect 9662 1710 9714 1762
rect 20862 1710 20914 1762
rect 21422 1710 21474 1762
<< metal2 >>
rect 672 49200 784 49800
rect 924 49308 1764 49364
rect 700 49140 756 49200
rect 924 49140 980 49308
rect 700 49084 980 49140
rect 1708 45332 1764 49308
rect 2016 49200 2128 49800
rect 4032 49200 4144 49800
rect 6048 49200 6160 49800
rect 7392 49200 7504 49800
rect 9408 49200 9520 49800
rect 11424 49200 11536 49800
rect 12768 49200 12880 49800
rect 14784 49200 14896 49800
rect 16128 49200 16240 49800
rect 18144 49200 18256 49800
rect 20160 49200 20272 49800
rect 21504 49200 21616 49800
rect 23520 49200 23632 49800
rect 25536 49200 25648 49800
rect 26880 49200 26992 49800
rect 28896 49200 29008 49800
rect 30912 49200 31024 49800
rect 32256 49200 32368 49800
rect 34272 49200 34384 49800
rect 35616 49200 35728 49800
rect 37632 49200 37744 49800
rect 39648 49200 39760 49800
rect 40992 49200 41104 49800
rect 43008 49200 43120 49800
rect 45024 49200 45136 49800
rect 46368 49200 46480 49800
rect 48384 49200 48496 49800
rect 49728 49200 49840 49800
rect 2044 45780 2100 49200
rect 3388 49140 3444 49150
rect 3388 47012 3444 49084
rect 2940 46956 3444 47012
rect 2268 45780 2324 45790
rect 2044 45778 2324 45780
rect 2044 45726 2270 45778
rect 2322 45726 2324 45778
rect 2044 45724 2324 45726
rect 2268 45714 2324 45724
rect 2492 45780 2548 45790
rect 1820 45668 1876 45678
rect 1820 45574 1876 45612
rect 1820 45332 1876 45342
rect 1708 45330 1876 45332
rect 1708 45278 1822 45330
rect 1874 45278 1876 45330
rect 1708 45276 1876 45278
rect 1820 45266 1876 45276
rect 2492 45330 2548 45724
rect 2940 45778 2996 46956
rect 2940 45726 2942 45778
rect 2994 45726 2996 45778
rect 2940 45714 2996 45726
rect 3052 46452 3108 46462
rect 2492 45278 2494 45330
rect 2546 45278 2548 45330
rect 2492 45266 2548 45278
rect 3052 44322 3108 46396
rect 4060 46002 4116 49200
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 6860 46116 6916 46126
rect 4060 45950 4062 46002
rect 4114 45950 4116 46002
rect 4060 45938 4116 45950
rect 5964 46004 6020 46014
rect 5964 46002 6132 46004
rect 5964 45950 5966 46002
rect 6018 45950 6132 46002
rect 5964 45948 6132 45950
rect 5964 45938 6020 45948
rect 4956 45892 5012 45902
rect 4956 45798 5012 45836
rect 3500 45668 3556 45678
rect 3164 45332 3220 45342
rect 3164 45238 3220 45276
rect 3500 45330 3556 45612
rect 4284 45668 4340 45678
rect 3500 45278 3502 45330
rect 3554 45278 3556 45330
rect 3500 45266 3556 45278
rect 4172 45556 4228 45566
rect 4060 44994 4116 45006
rect 4060 44942 4062 44994
rect 4114 44942 4116 44994
rect 3724 44436 3780 44446
rect 3724 44342 3780 44380
rect 3052 44270 3054 44322
rect 3106 44270 3108 44322
rect 2156 44210 2212 44222
rect 2156 44158 2158 44210
rect 2210 44158 2212 44210
rect 2156 43764 2212 44158
rect 2156 43698 2212 43708
rect 3052 43762 3108 44270
rect 4060 43876 4116 44942
rect 4172 44434 4228 45500
rect 4172 44382 4174 44434
rect 4226 44382 4228 44434
rect 4172 44370 4228 44382
rect 4284 45108 4340 45612
rect 4060 43810 4116 43820
rect 3052 43710 3054 43762
rect 3106 43710 3108 43762
rect 3052 43698 3108 43710
rect 4284 43762 4340 45052
rect 5516 45668 5572 45678
rect 5516 45330 5572 45612
rect 5516 45278 5518 45330
rect 5570 45278 5572 45330
rect 4508 44996 4564 45006
rect 4956 44996 5012 45006
rect 4508 44994 4900 44996
rect 4508 44942 4510 44994
rect 4562 44942 4900 44994
rect 4508 44940 4900 44942
rect 4508 44930 4564 44940
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4620 44100 4676 44110
rect 4620 44006 4676 44044
rect 4844 43988 4900 44940
rect 4956 44902 5012 44940
rect 5404 44994 5460 45006
rect 5404 44942 5406 44994
rect 5458 44942 5460 44994
rect 5068 44098 5124 44110
rect 5068 44046 5070 44098
rect 5122 44046 5124 44098
rect 5068 43988 5124 44046
rect 4844 43932 5012 43988
rect 4284 43710 4286 43762
rect 4338 43710 4340 43762
rect 3500 43428 3556 43438
rect 3500 43334 3556 43372
rect 3948 43426 4004 43438
rect 3948 43374 3950 43426
rect 4002 43374 4004 43426
rect 3948 42868 4004 43374
rect 3948 42802 4004 42812
rect 1820 42530 1876 42542
rect 1820 42478 1822 42530
rect 1874 42478 1876 42530
rect 1820 42420 1876 42478
rect 1820 42354 1876 42364
rect 4284 42196 4340 43710
rect 4844 43764 4900 43774
rect 4844 43670 4900 43708
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4508 42868 4564 42878
rect 4508 42774 4564 42812
rect 4284 42130 4340 42140
rect 4956 41636 5012 43932
rect 5068 43922 5124 43932
rect 5180 43876 5236 43886
rect 5180 43762 5236 43820
rect 5180 43710 5182 43762
rect 5234 43710 5236 43762
rect 5068 43652 5124 43662
rect 5068 42866 5124 43596
rect 5180 43540 5236 43710
rect 5180 43474 5236 43484
rect 5068 42814 5070 42866
rect 5122 42814 5124 42866
rect 5068 42802 5124 42814
rect 5404 43428 5460 44942
rect 5516 43764 5572 45278
rect 5740 45444 5796 45454
rect 5628 43764 5684 43774
rect 5516 43762 5684 43764
rect 5516 43710 5630 43762
rect 5682 43710 5684 43762
rect 5516 43708 5684 43710
rect 5628 43698 5684 43708
rect 5292 41858 5348 41870
rect 5292 41806 5294 41858
rect 5346 41806 5348 41858
rect 5292 41746 5348 41806
rect 5292 41694 5294 41746
rect 5346 41694 5348 41746
rect 5292 41682 5348 41694
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4956 41570 5012 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5404 39844 5460 43372
rect 5740 42866 5796 45388
rect 5740 42814 5742 42866
rect 5794 42814 5796 42866
rect 5740 42802 5796 42814
rect 5852 44324 5908 44334
rect 5852 44210 5908 44268
rect 5852 44158 5854 44210
rect 5906 44158 5908 44210
rect 5628 42196 5684 42206
rect 5628 41076 5684 42140
rect 5852 41746 5908 44158
rect 5852 41694 5854 41746
rect 5906 41694 5908 41746
rect 5852 41682 5908 41694
rect 5964 44098 6020 44110
rect 5964 44046 5966 44098
rect 6018 44046 6020 44098
rect 5628 41010 5684 41020
rect 5404 39778 5460 39788
rect 5964 39060 6020 44046
rect 6076 43652 6132 45948
rect 6860 45220 6916 46060
rect 6860 45218 7028 45220
rect 6860 45166 6862 45218
rect 6914 45166 7028 45218
rect 6860 45164 7028 45166
rect 6860 45154 6916 45164
rect 6188 45108 6244 45118
rect 6188 45014 6244 45052
rect 6524 44324 6580 44334
rect 6524 44230 6580 44268
rect 6748 43876 6804 43886
rect 6748 43762 6804 43820
rect 6748 43710 6750 43762
rect 6802 43710 6804 43762
rect 6748 43698 6804 43710
rect 6076 43586 6132 43596
rect 6188 43428 6244 43438
rect 6188 43426 6356 43428
rect 6188 43374 6190 43426
rect 6242 43374 6356 43426
rect 6188 43372 6356 43374
rect 6188 43362 6244 43372
rect 6188 42532 6244 42542
rect 6076 42530 6244 42532
rect 6076 42478 6190 42530
rect 6242 42478 6244 42530
rect 6076 42476 6244 42478
rect 6076 41748 6132 42476
rect 6188 42466 6244 42476
rect 6188 42196 6244 42206
rect 6188 41970 6244 42140
rect 6188 41918 6190 41970
rect 6242 41918 6244 41970
rect 6188 41906 6244 41918
rect 6300 41972 6356 43372
rect 6636 42980 6692 42990
rect 6636 42866 6692 42924
rect 6636 42814 6638 42866
rect 6690 42814 6692 42866
rect 6636 42802 6692 42814
rect 6300 41906 6356 41916
rect 6076 41682 6132 41692
rect 6636 41858 6692 41870
rect 6636 41806 6638 41858
rect 6690 41806 6692 41858
rect 5964 38994 6020 39004
rect 6412 41300 6468 41310
rect 1820 38946 1876 38958
rect 1820 38894 1822 38946
rect 1874 38894 1876 38946
rect 1820 38388 1876 38894
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 1820 38322 1876 38332
rect 6412 37940 6468 41244
rect 6636 40180 6692 41806
rect 6636 40114 6692 40124
rect 6748 41746 6804 41758
rect 6748 41694 6750 41746
rect 6802 41694 6804 41746
rect 6748 40962 6804 41694
rect 6748 40910 6750 40962
rect 6802 40910 6804 40962
rect 6748 38948 6804 40910
rect 6972 40178 7028 45164
rect 7308 44212 7364 44222
rect 7308 44118 7364 44156
rect 7420 43876 7476 49200
rect 7980 46004 8036 46014
rect 7420 43810 7476 43820
rect 7756 45220 7812 45230
rect 7308 43428 7364 43438
rect 7308 42868 7364 43372
rect 7308 42802 7364 42812
rect 7420 43314 7476 43326
rect 7420 43262 7422 43314
rect 7474 43262 7476 43314
rect 7084 42756 7140 42766
rect 7084 42662 7140 42700
rect 7420 42532 7476 43262
rect 7644 42868 7700 42878
rect 7196 42476 7476 42532
rect 7532 42530 7588 42542
rect 7532 42478 7534 42530
rect 7586 42478 7588 42530
rect 7084 41860 7140 41870
rect 7084 41766 7140 41804
rect 6972 40126 6974 40178
rect 7026 40126 7028 40178
rect 6972 40114 7028 40126
rect 7196 39396 7252 42476
rect 7532 42084 7588 42478
rect 7532 42018 7588 42028
rect 7420 41858 7476 41870
rect 7420 41806 7422 41858
rect 7474 41806 7476 41858
rect 7420 41748 7476 41806
rect 7308 41524 7364 41534
rect 7308 41298 7364 41468
rect 7420 41410 7476 41692
rect 7420 41358 7422 41410
rect 7474 41358 7476 41410
rect 7420 41346 7476 41358
rect 7308 41246 7310 41298
rect 7362 41246 7364 41298
rect 7308 41234 7364 41246
rect 7308 40628 7364 40638
rect 7644 40628 7700 42812
rect 7756 41298 7812 45164
rect 7868 44548 7924 44558
rect 7868 43764 7924 44492
rect 7868 41970 7924 43708
rect 7980 43650 8036 45948
rect 8764 45890 8820 45902
rect 8764 45838 8766 45890
rect 8818 45838 8820 45890
rect 8092 45780 8148 45790
rect 8092 45686 8148 45724
rect 8764 45108 8820 45838
rect 9436 45668 9492 49200
rect 11340 48244 11396 48254
rect 10668 48132 10724 48142
rect 9996 47796 10052 47806
rect 9996 45890 10052 47740
rect 9996 45838 9998 45890
rect 10050 45838 10052 45890
rect 9100 45612 9492 45668
rect 9548 45780 9604 45790
rect 8764 45042 8820 45052
rect 8988 45220 9044 45230
rect 8988 44994 9044 45164
rect 8988 44942 8990 44994
rect 9042 44942 9044 44994
rect 8988 44930 9044 44942
rect 8988 43764 9044 43774
rect 7980 43598 7982 43650
rect 8034 43598 8036 43650
rect 7980 42868 8036 43598
rect 8876 43652 8932 43662
rect 8876 43558 8932 43596
rect 8764 43540 8820 43550
rect 8540 43428 8596 43438
rect 8092 43316 8148 43326
rect 8540 43316 8596 43372
rect 8652 43316 8708 43326
rect 8092 43314 8260 43316
rect 8092 43262 8094 43314
rect 8146 43262 8260 43314
rect 8092 43260 8260 43262
rect 8092 43250 8148 43260
rect 7980 42802 8036 42812
rect 8204 42756 8260 43260
rect 8540 43314 8708 43316
rect 8540 43262 8654 43314
rect 8706 43262 8708 43314
rect 8540 43260 8708 43262
rect 7868 41918 7870 41970
rect 7922 41918 7924 41970
rect 7868 41746 7924 41918
rect 7868 41694 7870 41746
rect 7922 41694 7924 41746
rect 7868 41682 7924 41694
rect 7980 42642 8036 42654
rect 7980 42590 7982 42642
rect 8034 42590 8036 42642
rect 7756 41246 7758 41298
rect 7810 41246 7812 41298
rect 7756 41234 7812 41246
rect 7980 41412 8036 42590
rect 8092 42532 8148 42542
rect 8092 42438 8148 42476
rect 7308 40626 7700 40628
rect 7308 40574 7310 40626
rect 7362 40574 7700 40626
rect 7308 40572 7700 40574
rect 7756 40628 7812 40638
rect 7980 40628 8036 41356
rect 8092 41636 8148 41646
rect 8092 41298 8148 41580
rect 8204 41524 8260 42700
rect 8428 43092 8484 43102
rect 8316 41858 8372 41870
rect 8316 41806 8318 41858
rect 8370 41806 8372 41858
rect 8316 41746 8372 41806
rect 8316 41694 8318 41746
rect 8370 41694 8372 41746
rect 8316 41682 8372 41694
rect 8204 41468 8372 41524
rect 8092 41246 8094 41298
rect 8146 41246 8148 41298
rect 8092 41234 8148 41246
rect 7756 40626 8036 40628
rect 7756 40574 7758 40626
rect 7810 40574 8036 40626
rect 7756 40572 8036 40574
rect 7308 40562 7364 40572
rect 7756 40562 7812 40572
rect 8204 40404 8260 40414
rect 8204 40310 8260 40348
rect 8204 40178 8260 40190
rect 8204 40126 8206 40178
rect 8258 40126 8260 40178
rect 8204 39732 8260 40126
rect 8316 40068 8372 41468
rect 8428 41410 8484 43036
rect 8428 41358 8430 41410
rect 8482 41358 8484 41410
rect 8428 40178 8484 41358
rect 8428 40126 8430 40178
rect 8482 40126 8484 40178
rect 8428 40114 8484 40126
rect 8316 40002 8372 40012
rect 8316 39732 8372 39742
rect 8204 39730 8372 39732
rect 8204 39678 8318 39730
rect 8370 39678 8372 39730
rect 8204 39676 8372 39678
rect 8316 39666 8372 39676
rect 7196 39330 7252 39340
rect 6748 38882 6804 38892
rect 6412 37874 6468 37884
rect 1820 37378 1876 37390
rect 1820 37326 1822 37378
rect 1874 37326 1876 37378
rect 1820 37044 1876 37326
rect 8540 37268 8596 43260
rect 8652 43250 8708 43260
rect 8764 42978 8820 43484
rect 8876 43428 8932 43438
rect 8876 43334 8932 43372
rect 8764 42926 8766 42978
rect 8818 42926 8820 42978
rect 8764 42914 8820 42926
rect 8652 42644 8708 42654
rect 8652 42550 8708 42588
rect 8988 42420 9044 43708
rect 8876 42364 9044 42420
rect 8764 42196 8820 42206
rect 8652 41636 8708 41646
rect 8652 41298 8708 41580
rect 8652 41246 8654 41298
rect 8706 41246 8708 41298
rect 8652 41234 8708 41246
rect 8652 40628 8708 40638
rect 8764 40628 8820 42140
rect 8652 40626 8820 40628
rect 8652 40574 8654 40626
rect 8706 40574 8820 40626
rect 8652 40572 8820 40574
rect 8652 40562 8708 40572
rect 8764 39732 8820 39742
rect 8876 39732 8932 42364
rect 8988 42196 9044 42206
rect 9100 42196 9156 45612
rect 9548 44996 9604 45724
rect 9996 45332 10052 45838
rect 10668 45778 10724 48076
rect 10668 45726 10670 45778
rect 10722 45726 10724 45778
rect 10668 45556 10724 45726
rect 10668 45490 10724 45500
rect 10892 47684 10948 47694
rect 9436 44436 9492 44446
rect 8988 42194 9156 42196
rect 8988 42142 8990 42194
rect 9042 42142 9156 42194
rect 8988 42140 9156 42142
rect 9212 44434 9492 44436
rect 9212 44382 9438 44434
rect 9490 44382 9492 44434
rect 9212 44380 9492 44382
rect 8988 42130 9044 42140
rect 9100 41188 9156 41198
rect 9100 41094 9156 41132
rect 9100 40628 9156 40638
rect 9212 40628 9268 44380
rect 9436 44370 9492 44380
rect 9324 43092 9380 43102
rect 9324 42866 9380 43036
rect 9436 42980 9492 42990
rect 9548 42980 9604 44940
rect 9772 45106 9828 45118
rect 9772 45054 9774 45106
rect 9826 45054 9828 45106
rect 9660 44884 9716 44894
rect 9660 43764 9716 44828
rect 9660 43698 9716 43708
rect 9772 43540 9828 45054
rect 9996 44434 10052 45276
rect 10108 45108 10164 45118
rect 10108 45014 10164 45052
rect 10332 45106 10388 45118
rect 10332 45054 10334 45106
rect 10386 45054 10388 45106
rect 9996 44382 9998 44434
rect 10050 44382 10052 44434
rect 9996 44370 10052 44382
rect 10220 44994 10276 45006
rect 10220 44942 10222 44994
rect 10274 44942 10276 44994
rect 9884 43764 9940 43774
rect 10108 43764 10164 43774
rect 9884 43762 10108 43764
rect 9884 43710 9886 43762
rect 9938 43710 10108 43762
rect 9884 43708 10108 43710
rect 9884 43698 9940 43708
rect 9996 43540 10052 43550
rect 9436 42978 9604 42980
rect 9436 42926 9438 42978
rect 9490 42926 9604 42978
rect 9436 42924 9604 42926
rect 9660 43484 9828 43540
rect 9884 43538 10052 43540
rect 9884 43486 9998 43538
rect 10050 43486 10052 43538
rect 9884 43484 10052 43486
rect 9436 42914 9492 42924
rect 9324 42814 9326 42866
rect 9378 42814 9380 42866
rect 9324 42802 9380 42814
rect 9100 40626 9268 40628
rect 9100 40574 9102 40626
rect 9154 40574 9268 40626
rect 9100 40572 9268 40574
rect 9100 40562 9156 40572
rect 9212 40516 9268 40572
rect 9212 40450 9268 40460
rect 9436 42756 9492 42766
rect 8764 39730 8932 39732
rect 8764 39678 8766 39730
rect 8818 39678 8932 39730
rect 8764 39676 8932 39678
rect 9100 40178 9156 40190
rect 9100 40126 9102 40178
rect 9154 40126 9156 40178
rect 9100 39730 9156 40126
rect 9100 39678 9102 39730
rect 9154 39678 9156 39730
rect 8764 39666 8820 39676
rect 9100 39666 9156 39678
rect 9436 39172 9492 42700
rect 9660 42084 9716 43484
rect 9884 42756 9940 43484
rect 9996 43474 10052 43484
rect 9884 42690 9940 42700
rect 9996 42866 10052 42878
rect 9996 42814 9998 42866
rect 10050 42814 10052 42866
rect 9996 42644 10052 42814
rect 9996 42578 10052 42588
rect 9548 42028 9716 42084
rect 9996 42420 10052 42430
rect 9548 41524 9604 42028
rect 9660 41858 9716 41870
rect 9660 41806 9662 41858
rect 9714 41806 9716 41858
rect 9660 41748 9716 41806
rect 9996 41860 10052 42364
rect 9996 41794 10052 41804
rect 9660 41682 9716 41692
rect 9548 41468 9716 41524
rect 9548 41300 9604 41310
rect 9548 41206 9604 41244
rect 9660 40628 9716 41468
rect 9996 41186 10052 41198
rect 9996 41134 9998 41186
rect 10050 41134 10052 41186
rect 9996 41076 10052 41134
rect 9996 41010 10052 41020
rect 9660 40292 9716 40572
rect 10108 40404 10164 43708
rect 10220 42868 10276 44942
rect 10332 43764 10388 45054
rect 10332 43698 10388 43708
rect 10444 44324 10500 44334
rect 10220 42802 10276 42812
rect 10220 41972 10276 41982
rect 10220 41878 10276 41916
rect 10332 41972 10388 41982
rect 10444 41972 10500 44268
rect 10668 43988 10724 43998
rect 10556 43538 10612 43550
rect 10556 43486 10558 43538
rect 10610 43486 10612 43538
rect 10556 43092 10612 43486
rect 10556 43026 10612 43036
rect 10332 41970 10500 41972
rect 10332 41918 10334 41970
rect 10386 41918 10500 41970
rect 10332 41916 10500 41918
rect 10332 41524 10388 41916
rect 10332 41458 10388 41468
rect 10220 40628 10276 40638
rect 10220 40534 10276 40572
rect 10668 40626 10724 43932
rect 10780 42532 10836 42542
rect 10780 41298 10836 42476
rect 10892 42196 10948 47628
rect 11004 45106 11060 45118
rect 11004 45054 11006 45106
rect 11058 45054 11060 45106
rect 11004 44772 11060 45054
rect 11116 45108 11172 45118
rect 11116 45014 11172 45052
rect 11228 45106 11284 45118
rect 11228 45054 11230 45106
rect 11282 45054 11284 45106
rect 11004 44436 11060 44716
rect 11228 44548 11284 45054
rect 11228 44482 11284 44492
rect 11004 44370 11060 44380
rect 10892 42064 10948 42140
rect 11228 44212 11284 44222
rect 10780 41246 10782 41298
rect 10834 41246 10836 41298
rect 10780 41234 10836 41246
rect 10668 40574 10670 40626
rect 10722 40574 10724 40626
rect 10668 40562 10724 40574
rect 11228 40626 11284 44156
rect 11340 43650 11396 48188
rect 11452 47684 11508 49200
rect 11452 47618 11508 47628
rect 11900 47906 11956 47918
rect 11900 47854 11902 47906
rect 11954 47854 11956 47906
rect 11452 44996 11508 45006
rect 11452 44902 11508 44940
rect 11676 44884 11732 44894
rect 11676 44790 11732 44828
rect 11564 44548 11620 44558
rect 11452 44212 11508 44222
rect 11452 43988 11508 44156
rect 11452 43922 11508 43932
rect 11340 43598 11342 43650
rect 11394 43598 11396 43650
rect 11340 42980 11396 43598
rect 11340 42914 11396 42924
rect 11564 42980 11620 44492
rect 11564 42914 11620 42924
rect 11452 42532 11508 42542
rect 11340 42084 11396 42094
rect 11340 41524 11396 42028
rect 11340 41458 11396 41468
rect 11452 41858 11508 42476
rect 11452 41806 11454 41858
rect 11506 41806 11508 41858
rect 11452 41300 11508 41806
rect 11340 41244 11508 41300
rect 11564 42420 11620 42430
rect 11340 40964 11396 41244
rect 11340 40898 11396 40908
rect 11452 41076 11508 41086
rect 11228 40574 11230 40626
rect 11282 40574 11284 40626
rect 11228 40562 11284 40574
rect 11340 40516 11396 40526
rect 10108 40338 10164 40348
rect 10556 40404 10612 40414
rect 9884 40292 9940 40302
rect 9660 40290 9940 40292
rect 9660 40238 9886 40290
rect 9938 40238 9940 40290
rect 9660 40236 9940 40238
rect 9548 39732 9604 39742
rect 9548 39638 9604 39676
rect 9884 39508 9940 40236
rect 10556 40068 10612 40348
rect 10556 40012 10724 40068
rect 9996 39732 10052 39742
rect 10556 39732 10612 39742
rect 10052 39676 10164 39732
rect 9996 39600 10052 39676
rect 9884 39452 10052 39508
rect 9436 39106 9492 39116
rect 9996 39058 10052 39452
rect 9996 39006 9998 39058
rect 10050 39006 10052 39058
rect 9996 38994 10052 39006
rect 10108 38612 10164 39676
rect 10556 39638 10612 39676
rect 10108 38546 10164 38556
rect 10444 39172 10500 39182
rect 10444 39058 10500 39116
rect 10444 39006 10446 39058
rect 10498 39006 10500 39058
rect 10444 37380 10500 39006
rect 10556 38164 10612 38174
rect 10668 38164 10724 40012
rect 11340 39508 11396 40460
rect 11452 39730 11508 41020
rect 11452 39678 11454 39730
rect 11506 39678 11508 39730
rect 11452 39666 11508 39678
rect 11340 39452 11508 39508
rect 11004 39396 11060 39406
rect 11004 39394 11172 39396
rect 11004 39342 11006 39394
rect 11058 39342 11172 39394
rect 11004 39340 11172 39342
rect 11004 39330 11060 39340
rect 10892 38722 10948 38734
rect 10892 38670 10894 38722
rect 10946 38670 10948 38722
rect 10892 38612 10948 38670
rect 10892 38546 10948 38556
rect 11004 38610 11060 38622
rect 11004 38558 11006 38610
rect 11058 38558 11060 38610
rect 10612 38108 10724 38164
rect 11004 38162 11060 38558
rect 11004 38110 11006 38162
rect 11058 38110 11060 38162
rect 10556 38070 10612 38108
rect 11004 38098 11060 38110
rect 10444 37314 10500 37324
rect 8540 37202 8596 37212
rect 1820 36978 1876 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 11116 36820 11172 39340
rect 11340 39060 11396 39070
rect 11340 38966 11396 39004
rect 11452 37492 11508 39452
rect 11564 37716 11620 42364
rect 11900 41636 11956 47854
rect 12796 47906 12852 49200
rect 16716 48020 16772 48030
rect 12796 47854 12798 47906
rect 12850 47854 12852 47906
rect 12796 47842 12852 47854
rect 14028 47908 14084 47918
rect 12796 46564 12852 46574
rect 12236 46452 12292 46462
rect 12124 45780 12180 45790
rect 12124 45444 12180 45724
rect 12124 44434 12180 45388
rect 12236 45330 12292 46396
rect 12796 46002 12852 46508
rect 12796 45950 12798 46002
rect 12850 45950 12852 46002
rect 12796 45938 12852 45950
rect 13580 45892 13636 45902
rect 13580 45798 13636 45836
rect 12236 45278 12238 45330
rect 12290 45278 12292 45330
rect 12236 45266 12292 45278
rect 12124 44382 12126 44434
rect 12178 44382 12180 44434
rect 12124 44370 12180 44382
rect 12908 44324 12964 44334
rect 12908 44322 13076 44324
rect 12908 44270 12910 44322
rect 12962 44270 13076 44322
rect 12908 44268 13076 44270
rect 12908 44258 12964 44268
rect 12572 43428 12628 43438
rect 12124 42642 12180 42654
rect 12124 42590 12126 42642
rect 12178 42590 12180 42642
rect 12124 42420 12180 42590
rect 12124 42354 12180 42364
rect 12572 42084 12628 43372
rect 12908 42754 12964 42766
rect 12908 42702 12910 42754
rect 12962 42702 12964 42754
rect 12908 42532 12964 42702
rect 12908 42466 12964 42476
rect 12012 41860 12068 41870
rect 12012 41858 12516 41860
rect 12012 41806 12014 41858
rect 12066 41806 12516 41858
rect 12012 41804 12516 41806
rect 12012 41794 12068 41804
rect 11900 41580 12068 41636
rect 11676 41188 11732 41198
rect 11676 38610 11732 41132
rect 11900 40292 11956 40302
rect 11676 38558 11678 38610
rect 11730 38558 11732 38610
rect 11676 38546 11732 38558
rect 11788 40290 11956 40292
rect 11788 40238 11902 40290
rect 11954 40238 11956 40290
rect 11788 40236 11956 40238
rect 11564 37650 11620 37660
rect 11452 37426 11508 37436
rect 11116 36754 11172 36764
rect 5852 36148 5908 36158
rect 1820 35810 1876 35822
rect 1820 35758 1822 35810
rect 1874 35758 1876 35810
rect 1820 35028 1876 35758
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1820 34962 1876 34972
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1820 33122 1876 33134
rect 1820 33070 1822 33122
rect 1874 33070 1876 33122
rect 1820 33012 1876 33070
rect 1820 32946 1876 32956
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1820 29986 1876 29998
rect 1820 29934 1822 29986
rect 1874 29934 1876 29986
rect 1820 29652 1876 29934
rect 1820 29586 1876 29596
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 1820 28418 1876 28430
rect 1820 28366 1822 28418
rect 1874 28366 1876 28418
rect 1820 28308 1876 28366
rect 1820 28242 1876 28252
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 1820 26850 1876 26862
rect 1820 26798 1822 26850
rect 1874 26798 1876 26850
rect 1820 26292 1876 26798
rect 1820 26226 1876 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1820 24834 1876 24846
rect 1820 24782 1822 24834
rect 1874 24782 1876 24834
rect 1820 24276 1876 24782
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 1820 24210 1876 24220
rect 3052 23380 3108 23390
rect 3052 23154 3108 23324
rect 3500 23380 3556 23390
rect 3500 23286 3556 23324
rect 3052 23102 3054 23154
rect 3106 23102 3108 23154
rect 3052 23090 3108 23102
rect 2044 23042 2100 23054
rect 2044 22990 2046 23042
rect 2098 22990 2100 23042
rect 2044 22932 2100 22990
rect 2044 22866 2100 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1820 21698 1876 21710
rect 1820 21646 1822 21698
rect 1874 21646 1876 21698
rect 1820 20916 1876 21646
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 1820 20850 1876 20860
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 1820 19010 1876 19022
rect 1820 18958 1822 19010
rect 1874 18958 1876 19010
rect 1820 18900 1876 18958
rect 1820 18834 1876 18844
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1820 17556 1876 17566
rect 1820 17462 1876 17500
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1820 15874 1876 15886
rect 1820 15822 1822 15874
rect 1874 15822 1876 15874
rect 1820 15540 1876 15822
rect 1820 15474 1876 15484
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 1820 14306 1876 14318
rect 1820 14254 1822 14306
rect 1874 14254 1876 14306
rect 1820 14196 1876 14254
rect 1820 14130 1876 14140
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 1820 10722 1876 10734
rect 1820 10670 1822 10722
rect 1874 10670 1876 10722
rect 1820 10164 1876 10670
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 1820 10098 1876 10108
rect 1820 9154 1876 9166
rect 1820 9102 1822 9154
rect 1874 9102 1876 9154
rect 1820 8820 1876 9102
rect 1820 8754 1876 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 1820 7586 1876 7598
rect 1820 7534 1822 7586
rect 1874 7534 1876 7586
rect 1820 6804 1876 7534
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 1820 6738 1876 6748
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 1820 4450 1876 4462
rect 1820 4398 1822 4450
rect 1874 4398 1876 4450
rect 1372 3556 1428 3566
rect 28 2324 84 2334
rect 28 800 84 2268
rect 1372 800 1428 3500
rect 1820 3444 1876 4398
rect 2492 4450 2548 4462
rect 2492 4398 2494 4450
rect 2546 4398 2548 4450
rect 2156 3556 2212 3566
rect 2156 3462 2212 3500
rect 1820 3378 1876 3388
rect 2492 2324 2548 4398
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 3052 3668 3108 3678
rect 3052 3554 3108 3612
rect 4284 3668 4340 3678
rect 4284 3574 4340 3612
rect 5852 3668 5908 36092
rect 11228 35588 11284 35598
rect 11228 23380 11284 35532
rect 11788 35588 11844 40236
rect 11900 40226 11956 40236
rect 11900 39956 11956 39966
rect 11900 39058 11956 39900
rect 12012 39506 12068 41580
rect 12012 39454 12014 39506
rect 12066 39454 12068 39506
rect 12012 39442 12068 39454
rect 12124 40404 12180 40414
rect 12124 39284 12180 40348
rect 11900 39006 11902 39058
rect 11954 39006 11956 39058
rect 11900 38994 11956 39006
rect 12012 39228 12180 39284
rect 12348 40068 12404 40078
rect 12012 38612 12068 39228
rect 12348 39058 12404 40012
rect 12348 39006 12350 39058
rect 12402 39006 12404 39058
rect 12348 38994 12404 39006
rect 12460 38668 12516 41804
rect 12572 39956 12628 42028
rect 12908 41412 12964 41422
rect 12908 41298 12964 41356
rect 12908 41246 12910 41298
rect 12962 41246 12964 41298
rect 12908 41234 12964 41246
rect 13020 40180 13076 44268
rect 13692 44210 13748 44222
rect 13692 44158 13694 44210
rect 13746 44158 13748 44210
rect 13692 43540 13748 44158
rect 13916 44100 13972 44110
rect 13468 43428 13524 43438
rect 13468 43334 13524 43372
rect 13692 43204 13748 43484
rect 13692 43138 13748 43148
rect 13804 44098 13972 44100
rect 13804 44046 13918 44098
rect 13970 44046 13972 44098
rect 13804 44044 13972 44046
rect 13804 42980 13860 44044
rect 13916 44034 13972 44044
rect 14028 43764 14084 47852
rect 15708 47572 15764 47582
rect 14476 45892 14532 45902
rect 14252 44546 14308 44558
rect 14252 44494 14254 44546
rect 14306 44494 14308 44546
rect 14140 44100 14196 44110
rect 14140 44006 14196 44044
rect 14028 43708 14196 43764
rect 14028 43540 14084 43550
rect 14028 43426 14084 43484
rect 14028 43374 14030 43426
rect 14082 43374 14084 43426
rect 14028 43362 14084 43374
rect 13692 42924 13860 42980
rect 13916 42980 13972 42990
rect 13692 41748 13748 42924
rect 13916 42420 13972 42924
rect 14140 42868 14196 43708
rect 13916 42354 13972 42364
rect 14028 42866 14196 42868
rect 14028 42814 14142 42866
rect 14194 42814 14196 42866
rect 14028 42812 14196 42814
rect 13020 40114 13076 40124
rect 13244 41412 13300 41422
rect 12572 39890 12628 39900
rect 12796 39620 12852 39630
rect 12572 39396 12628 39406
rect 12572 39394 12740 39396
rect 12572 39342 12574 39394
rect 12626 39342 12740 39394
rect 12572 39340 12740 39342
rect 12572 39330 12628 39340
rect 12012 38162 12068 38556
rect 12012 38110 12014 38162
rect 12066 38110 12068 38162
rect 12012 38098 12068 38110
rect 12124 38612 12516 38668
rect 12124 36148 12180 38612
rect 12572 38274 12628 38286
rect 12572 38222 12574 38274
rect 12626 38222 12628 38274
rect 12572 38162 12628 38222
rect 12572 38110 12574 38162
rect 12626 38110 12628 38162
rect 12572 38098 12628 38110
rect 12684 38164 12740 39340
rect 12796 39058 12852 39564
rect 12796 39006 12798 39058
rect 12850 39006 12852 39058
rect 12796 38994 12852 39006
rect 12908 39508 12964 39518
rect 12684 37156 12740 38108
rect 12908 37492 12964 39452
rect 13244 38834 13300 41356
rect 13692 41188 13748 41692
rect 13692 41122 13748 41132
rect 13804 42308 13860 42318
rect 13804 41074 13860 42252
rect 13804 41022 13806 41074
rect 13858 41022 13860 41074
rect 13804 41010 13860 41022
rect 13692 40516 13748 40526
rect 13692 39730 13748 40460
rect 13692 39678 13694 39730
rect 13746 39678 13748 39730
rect 13692 39666 13748 39678
rect 14028 39732 14084 42812
rect 14140 42802 14196 42812
rect 14252 41186 14308 44494
rect 14364 44210 14420 44222
rect 14364 44158 14366 44210
rect 14418 44158 14420 44210
rect 14364 43092 14420 44158
rect 14364 43026 14420 43036
rect 14476 42866 14532 45836
rect 14924 45332 14980 45342
rect 14588 45108 14644 45118
rect 14588 45014 14644 45052
rect 14476 42814 14478 42866
rect 14530 42814 14532 42866
rect 14476 42802 14532 42814
rect 14588 44884 14644 44894
rect 14364 42756 14420 42766
rect 14364 42662 14420 42700
rect 14588 42530 14644 44828
rect 14588 42478 14590 42530
rect 14642 42478 14644 42530
rect 14252 41134 14254 41186
rect 14306 41134 14308 41186
rect 14252 41122 14308 41134
rect 14364 42196 14420 42206
rect 14364 41188 14420 42140
rect 14476 41970 14532 41982
rect 14476 41918 14478 41970
rect 14530 41918 14532 41970
rect 14476 41748 14532 41918
rect 14588 41860 14644 42478
rect 14588 41794 14644 41804
rect 14924 42532 14980 45276
rect 15372 45332 15428 45342
rect 15372 45106 15428 45276
rect 15372 45054 15374 45106
rect 15426 45054 15428 45106
rect 15372 45042 15428 45054
rect 15148 44436 15204 44446
rect 14924 41970 14980 42476
rect 14924 41918 14926 41970
rect 14978 41918 14980 41970
rect 14476 41682 14532 41692
rect 14924 41412 14980 41918
rect 14924 41346 14980 41356
rect 15036 42644 15092 42654
rect 14700 41188 14756 41198
rect 14364 41186 14756 41188
rect 14364 41134 14702 41186
rect 14754 41134 14756 41186
rect 14364 41132 14756 41134
rect 14028 39666 14084 39676
rect 14140 40964 14196 40974
rect 14140 39618 14196 40908
rect 14364 40628 14420 41132
rect 14700 41122 14756 41132
rect 14812 40962 14868 40974
rect 14812 40910 14814 40962
rect 14866 40910 14868 40962
rect 14812 40852 14868 40910
rect 14924 40964 14980 40974
rect 14924 40870 14980 40908
rect 14812 40786 14868 40796
rect 14252 40402 14308 40414
rect 14252 40350 14254 40402
rect 14306 40350 14308 40402
rect 14252 39730 14308 40350
rect 14364 40292 14420 40572
rect 14924 40404 14980 40414
rect 14924 40310 14980 40348
rect 14364 40226 14420 40236
rect 14252 39678 14254 39730
rect 14306 39678 14308 39730
rect 14252 39666 14308 39678
rect 15036 39732 15092 42588
rect 15148 41636 15204 44380
rect 15596 44436 15652 44446
rect 15596 44322 15652 44380
rect 15596 44270 15598 44322
rect 15650 44270 15652 44322
rect 15596 44258 15652 44270
rect 15708 43540 15764 47516
rect 16604 47460 16660 47470
rect 16044 47348 16100 47358
rect 15932 45892 15988 45902
rect 15932 45798 15988 45836
rect 15820 45220 15876 45230
rect 15820 44434 15876 45164
rect 15932 44996 15988 45006
rect 15932 44902 15988 44940
rect 15820 44382 15822 44434
rect 15874 44382 15876 44434
rect 15820 44370 15876 44382
rect 15932 44322 15988 44334
rect 15932 44270 15934 44322
rect 15986 44270 15988 44322
rect 15596 43484 15764 43540
rect 15820 44212 15876 44222
rect 15260 42980 15316 42990
rect 15260 42754 15316 42924
rect 15260 42702 15262 42754
rect 15314 42702 15316 42754
rect 15260 42690 15316 42702
rect 15148 41570 15204 41580
rect 15372 42530 15428 42542
rect 15372 42478 15374 42530
rect 15426 42478 15428 42530
rect 15036 39666 15092 39676
rect 15148 41412 15204 41422
rect 14140 39566 14142 39618
rect 14194 39566 14196 39618
rect 14028 39060 14084 39070
rect 14028 38946 14084 39004
rect 14028 38894 14030 38946
rect 14082 38894 14084 38946
rect 14028 38882 14084 38894
rect 13244 38782 13246 38834
rect 13298 38782 13300 38834
rect 13244 38668 13300 38782
rect 13132 38612 13300 38668
rect 13132 38274 13188 38612
rect 13132 38222 13134 38274
rect 13186 38222 13188 38274
rect 13132 38210 13188 38222
rect 13020 38164 13076 38174
rect 13020 38070 13076 38108
rect 13916 37826 13972 37838
rect 13916 37774 13918 37826
rect 13970 37774 13972 37826
rect 13132 37492 13188 37502
rect 12908 37490 13188 37492
rect 12908 37438 13134 37490
rect 13186 37438 13188 37490
rect 12908 37436 13188 37438
rect 13132 37426 13188 37436
rect 12684 37090 12740 37100
rect 13692 37154 13748 37166
rect 13692 37102 13694 37154
rect 13746 37102 13748 37154
rect 13692 36260 13748 37102
rect 13916 36596 13972 37774
rect 14140 37490 14196 39566
rect 14812 39618 14868 39630
rect 14812 39566 14814 39618
rect 14866 39566 14868 39618
rect 14140 37438 14142 37490
rect 14194 37438 14196 37490
rect 14140 37426 14196 37438
rect 14252 39396 14308 39406
rect 14252 38836 14308 39340
rect 14252 38162 14308 38780
rect 14252 38110 14254 38162
rect 14306 38110 14308 38162
rect 14252 37042 14308 38110
rect 14252 36990 14254 37042
rect 14306 36990 14308 37042
rect 14252 36978 14308 36990
rect 14364 39394 14420 39406
rect 14364 39342 14366 39394
rect 14418 39342 14420 39394
rect 14364 36708 14420 39342
rect 14812 39172 14868 39566
rect 15148 39620 15204 41356
rect 15372 40404 15428 42478
rect 15484 42530 15540 42542
rect 15484 42478 15486 42530
rect 15538 42478 15540 42530
rect 15484 42196 15540 42478
rect 15484 42130 15540 42140
rect 15596 41860 15652 43484
rect 15708 43316 15764 43326
rect 15708 43092 15764 43260
rect 15708 43026 15764 43036
rect 15708 42868 15764 42878
rect 15708 42754 15764 42812
rect 15708 42702 15710 42754
rect 15762 42702 15764 42754
rect 15708 42690 15764 42702
rect 15820 42084 15876 44156
rect 15484 41804 15652 41860
rect 15708 42028 15876 42084
rect 15484 41410 15540 41804
rect 15484 41358 15486 41410
rect 15538 41358 15540 41410
rect 15484 41076 15540 41358
rect 15596 41636 15652 41646
rect 15596 41410 15652 41580
rect 15596 41358 15598 41410
rect 15650 41358 15652 41410
rect 15596 41346 15652 41358
rect 15484 41010 15540 41020
rect 15484 40628 15540 40638
rect 15708 40628 15764 42028
rect 15820 41860 15876 41870
rect 15820 41410 15876 41804
rect 15820 41358 15822 41410
rect 15874 41358 15876 41410
rect 15820 41188 15876 41358
rect 15932 41412 15988 44270
rect 16044 43652 16100 47292
rect 16268 46228 16324 46238
rect 16268 44996 16324 46172
rect 16492 45890 16548 45902
rect 16492 45838 16494 45890
rect 16546 45838 16548 45890
rect 16156 44994 16324 44996
rect 16156 44942 16270 44994
rect 16322 44942 16324 44994
rect 16380 45668 16436 45678
rect 16380 45108 16436 45612
rect 16492 45332 16548 45838
rect 16492 45266 16548 45276
rect 16380 44976 16436 45052
rect 16156 44940 16324 44942
rect 16156 44212 16212 44940
rect 16268 44930 16324 44940
rect 16156 44146 16212 44156
rect 16492 44772 16548 44782
rect 16268 44100 16324 44110
rect 16268 44006 16324 44044
rect 16044 43596 16324 43652
rect 16156 43426 16212 43438
rect 16156 43374 16158 43426
rect 16210 43374 16212 43426
rect 16156 43092 16212 43374
rect 16156 43026 16212 43036
rect 16044 42868 16100 42878
rect 16044 42754 16100 42812
rect 16044 42702 16046 42754
rect 16098 42702 16100 42754
rect 16044 42420 16100 42702
rect 16044 42354 16100 42364
rect 16268 42084 16324 43596
rect 16156 41636 16212 41646
rect 15932 41356 16100 41412
rect 15820 41122 15876 41132
rect 15932 41186 15988 41198
rect 15932 41134 15934 41186
rect 15986 41134 15988 41186
rect 15484 40626 15708 40628
rect 15484 40574 15486 40626
rect 15538 40574 15708 40626
rect 15484 40572 15708 40574
rect 15484 40562 15540 40572
rect 15708 40496 15764 40572
rect 15820 40740 15876 40750
rect 15820 40514 15876 40684
rect 15820 40462 15822 40514
rect 15874 40462 15876 40514
rect 15820 40450 15876 40462
rect 15372 40348 15540 40404
rect 15148 39508 15204 39564
rect 15372 40180 15428 40190
rect 15260 39508 15316 39518
rect 15148 39506 15316 39508
rect 15148 39454 15262 39506
rect 15314 39454 15316 39506
rect 15148 39452 15316 39454
rect 15260 39442 15316 39452
rect 14812 39106 14868 39116
rect 14812 37940 14868 37950
rect 14812 37846 14868 37884
rect 14924 37940 14980 37950
rect 14924 37938 15092 37940
rect 14924 37886 14926 37938
rect 14978 37886 15092 37938
rect 14924 37884 15092 37886
rect 14924 37874 14980 37884
rect 14588 37492 14644 37502
rect 14588 37398 14644 37436
rect 14924 37156 14980 37166
rect 14924 37062 14980 37100
rect 14364 36642 14420 36652
rect 14700 37042 14756 37054
rect 14700 36990 14702 37042
rect 14754 36990 14756 37042
rect 13916 36530 13972 36540
rect 14700 36594 14756 36990
rect 14700 36542 14702 36594
rect 14754 36542 14756 36594
rect 13692 36194 13748 36204
rect 12124 36082 12180 36092
rect 14700 36036 14756 36542
rect 15036 36596 15092 37884
rect 15260 36932 15316 36942
rect 15260 36708 15316 36876
rect 15260 36642 15316 36652
rect 15372 36596 15428 40124
rect 15484 39172 15540 40348
rect 15820 40180 15876 40190
rect 15596 40068 15652 40078
rect 15596 39732 15652 40012
rect 15596 39618 15652 39676
rect 15596 39566 15598 39618
rect 15650 39566 15652 39618
rect 15596 39554 15652 39566
rect 15708 39956 15764 39966
rect 15708 39730 15764 39900
rect 15708 39678 15710 39730
rect 15762 39678 15764 39730
rect 15484 39106 15540 39116
rect 15596 39284 15652 39294
rect 15596 38164 15652 39228
rect 15596 38098 15652 38108
rect 15484 38050 15540 38062
rect 15484 37998 15486 38050
rect 15538 37998 15540 38050
rect 15484 37492 15540 37998
rect 15484 37426 15540 37436
rect 15484 37268 15540 37278
rect 15484 37174 15540 37212
rect 15596 36596 15652 36606
rect 15372 36594 15652 36596
rect 15372 36542 15598 36594
rect 15650 36542 15652 36594
rect 15372 36540 15652 36542
rect 15036 36530 15092 36540
rect 15148 36484 15204 36494
rect 15148 36260 15204 36428
rect 15596 36484 15652 36540
rect 15596 36418 15652 36428
rect 15148 36258 15316 36260
rect 15148 36206 15150 36258
rect 15202 36206 15316 36258
rect 15148 36204 15316 36206
rect 15148 36194 15204 36204
rect 14700 35970 14756 35980
rect 15260 36036 15316 36204
rect 15260 35970 15316 35980
rect 11788 35522 11844 35532
rect 15708 35252 15764 39678
rect 15820 39618 15876 40124
rect 15820 39566 15822 39618
rect 15874 39566 15876 39618
rect 15820 39554 15876 39566
rect 15820 39396 15876 39406
rect 15820 35924 15876 39340
rect 15932 37716 15988 41134
rect 16044 39060 16100 41356
rect 16156 41188 16212 41580
rect 16156 39284 16212 41132
rect 16268 40740 16324 42028
rect 16380 41970 16436 41982
rect 16380 41918 16382 41970
rect 16434 41918 16436 41970
rect 16380 41860 16436 41918
rect 16380 41794 16436 41804
rect 16380 41636 16436 41646
rect 16380 41412 16436 41580
rect 16380 41346 16436 41356
rect 16268 40674 16324 40684
rect 16380 41076 16436 41086
rect 16380 40514 16436 41020
rect 16492 40626 16548 44716
rect 16604 43540 16660 47404
rect 16716 45220 16772 47964
rect 17836 45780 17892 45790
rect 17500 45668 17556 45678
rect 17500 45574 17556 45612
rect 16716 45154 16772 45164
rect 17724 45106 17780 45118
rect 17724 45054 17726 45106
rect 17778 45054 17780 45106
rect 16828 44324 16884 44334
rect 16828 43764 16884 44268
rect 16828 43698 16884 43708
rect 17388 44212 17444 44222
rect 16604 43484 16772 43540
rect 16604 43316 16660 43326
rect 16604 42866 16660 43260
rect 16604 42814 16606 42866
rect 16658 42814 16660 42866
rect 16604 42532 16660 42814
rect 16604 42466 16660 42476
rect 16716 41970 16772 43484
rect 16716 41918 16718 41970
rect 16770 41918 16772 41970
rect 16604 41524 16660 41534
rect 16604 41298 16660 41468
rect 16604 41246 16606 41298
rect 16658 41246 16660 41298
rect 16604 41234 16660 41246
rect 16716 41300 16772 41918
rect 16716 41234 16772 41244
rect 16828 43538 16884 43550
rect 16828 43486 16830 43538
rect 16882 43486 16884 43538
rect 16828 43316 16884 43486
rect 16828 42084 16884 43260
rect 16492 40574 16494 40626
rect 16546 40574 16548 40626
rect 16492 40562 16548 40574
rect 16604 40628 16660 40638
rect 16380 40462 16382 40514
rect 16434 40462 16436 40514
rect 16380 40450 16436 40462
rect 16604 40402 16660 40572
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 16604 40338 16660 40350
rect 16380 39618 16436 39630
rect 16380 39566 16382 39618
rect 16434 39566 16436 39618
rect 16380 39508 16436 39566
rect 16380 39442 16436 39452
rect 16828 39396 16884 42028
rect 16940 41858 16996 41870
rect 16940 41806 16942 41858
rect 16994 41806 16996 41858
rect 16940 40740 16996 41806
rect 16940 40674 16996 40684
rect 17052 41860 17108 41870
rect 16940 40516 16996 40526
rect 16940 40422 16996 40460
rect 17052 40180 17108 41804
rect 16828 39330 16884 39340
rect 16940 40124 17108 40180
rect 16156 39218 16212 39228
rect 16044 38836 16100 39004
rect 16716 39060 16772 39070
rect 16044 38770 16100 38780
rect 16156 38948 16212 38958
rect 16156 38722 16212 38892
rect 16716 38946 16772 39004
rect 16716 38894 16718 38946
rect 16770 38894 16772 38946
rect 16716 38882 16772 38894
rect 16828 38946 16884 38958
rect 16828 38894 16830 38946
rect 16882 38894 16884 38946
rect 16156 38670 16158 38722
rect 16210 38670 16212 38722
rect 16156 38658 16212 38670
rect 16716 38052 16772 38062
rect 16268 37940 16324 37950
rect 16268 37938 16548 37940
rect 16268 37886 16270 37938
rect 16322 37886 16548 37938
rect 16268 37884 16548 37886
rect 16268 37874 16324 37884
rect 15932 37660 16436 37716
rect 15932 37156 15988 37166
rect 15932 36932 15988 37100
rect 16044 37044 16100 37054
rect 16044 36950 16100 36988
rect 15932 36866 15988 36876
rect 16156 36708 16212 36718
rect 16156 36594 16212 36652
rect 16156 36542 16158 36594
rect 16210 36542 16212 36594
rect 16156 36530 16212 36542
rect 16156 35924 16212 35934
rect 15820 35922 16212 35924
rect 15820 35870 16158 35922
rect 16210 35870 16212 35922
rect 15820 35868 16212 35870
rect 16380 35924 16436 37660
rect 16492 36708 16548 37884
rect 16604 37268 16660 37278
rect 16604 37174 16660 37212
rect 16716 37044 16772 37996
rect 16716 36978 16772 36988
rect 16604 36708 16660 36718
rect 16492 36706 16660 36708
rect 16492 36654 16606 36706
rect 16658 36654 16660 36706
rect 16492 36652 16660 36654
rect 16604 36642 16660 36652
rect 16828 36708 16884 38894
rect 16828 36642 16884 36652
rect 16940 37378 16996 40124
rect 17388 39956 17444 44156
rect 17388 39890 17444 39900
rect 17500 44210 17556 44222
rect 17500 44158 17502 44210
rect 17554 44158 17556 44210
rect 17276 39844 17332 39854
rect 17164 39620 17220 39630
rect 17164 39526 17220 39564
rect 17052 38836 17108 38846
rect 17052 38742 17108 38780
rect 16940 37326 16942 37378
rect 16994 37326 16996 37378
rect 16716 36484 16772 36494
rect 16772 36428 16884 36484
rect 16716 36390 16772 36428
rect 16604 35924 16660 35934
rect 16380 35922 16660 35924
rect 16380 35870 16606 35922
rect 16658 35870 16660 35922
rect 16380 35868 16660 35870
rect 16156 35858 16212 35868
rect 16604 35700 16660 35868
rect 16828 35812 16884 36428
rect 16940 35924 16996 37326
rect 17276 38164 17332 39788
rect 17388 39732 17444 39742
rect 17500 39732 17556 44158
rect 17724 43204 17780 45054
rect 17724 43138 17780 43148
rect 17836 43538 17892 45724
rect 18172 45332 18228 49200
rect 19404 46788 19460 46798
rect 18956 45668 19012 45678
rect 18060 45276 18228 45332
rect 18396 45444 18452 45454
rect 17836 43486 17838 43538
rect 17890 43486 17892 43538
rect 17724 42084 17780 42094
rect 17724 41858 17780 42028
rect 17724 41806 17726 41858
rect 17778 41806 17780 41858
rect 17724 41794 17780 41806
rect 17836 41524 17892 43486
rect 17948 45106 18004 45118
rect 17948 45054 17950 45106
rect 18002 45054 18004 45106
rect 17948 41860 18004 45054
rect 18060 42308 18116 45276
rect 18396 45220 18452 45388
rect 18172 45106 18228 45118
rect 18172 45054 18174 45106
rect 18226 45054 18228 45106
rect 18396 45088 18452 45164
rect 18956 45106 19012 45612
rect 18172 43988 18228 45054
rect 18956 45054 18958 45106
rect 19010 45054 19012 45106
rect 18956 45042 19012 45054
rect 18172 43922 18228 43932
rect 18284 44882 18340 44894
rect 18284 44830 18286 44882
rect 18338 44830 18340 44882
rect 18060 42242 18116 42252
rect 18172 43204 18228 43214
rect 17948 41794 18004 41804
rect 17836 41458 17892 41468
rect 18060 41748 18116 41758
rect 17724 41412 17780 41422
rect 17724 40290 17780 41356
rect 17724 40238 17726 40290
rect 17778 40238 17780 40290
rect 17724 40226 17780 40238
rect 17948 40292 18004 40302
rect 17444 39676 17556 39732
rect 17388 39666 17444 39676
rect 17276 36482 17332 38108
rect 17500 39508 17556 39518
rect 17500 37044 17556 39452
rect 17948 39508 18004 40236
rect 17612 39172 17668 39182
rect 17612 37266 17668 39116
rect 17948 39058 18004 39452
rect 17948 39006 17950 39058
rect 18002 39006 18004 39058
rect 17836 38948 17892 38958
rect 17836 38854 17892 38892
rect 17724 38836 17780 38846
rect 17724 38742 17780 38780
rect 17948 37828 18004 39006
rect 17948 37762 18004 37772
rect 18060 37492 18116 41692
rect 18172 40404 18228 43148
rect 18284 42084 18340 44830
rect 19180 43988 19236 43998
rect 18284 42018 18340 42028
rect 18508 43426 18564 43438
rect 18508 43374 18510 43426
rect 18562 43374 18564 43426
rect 18508 41972 18564 43374
rect 18508 41906 18564 41916
rect 18620 42868 18676 42878
rect 18172 40338 18228 40348
rect 18508 39956 18564 39966
rect 18396 39396 18452 39406
rect 18396 38834 18452 39340
rect 18396 38782 18398 38834
rect 18450 38782 18452 38834
rect 18396 38770 18452 38782
rect 18508 38724 18564 39900
rect 18508 38658 18564 38668
rect 18620 38668 18676 42812
rect 18732 42642 18788 42654
rect 18732 42590 18734 42642
rect 18786 42590 18788 42642
rect 18732 41860 18788 42590
rect 19068 41860 19124 41870
rect 18732 41804 19068 41860
rect 18732 41300 18788 41310
rect 18732 41206 18788 41244
rect 18956 40180 19012 40190
rect 18956 39058 19012 40124
rect 18956 39006 18958 39058
rect 19010 39006 19012 39058
rect 18956 38994 19012 39006
rect 19068 39058 19124 41804
rect 19068 39006 19070 39058
rect 19122 39006 19124 39058
rect 19068 38994 19124 39006
rect 18844 38836 18900 38874
rect 18844 38770 18900 38780
rect 19180 38836 19236 43932
rect 19292 39844 19348 39854
rect 19292 39730 19348 39788
rect 19292 39678 19294 39730
rect 19346 39678 19348 39730
rect 19292 39666 19348 39678
rect 19292 39060 19348 39070
rect 19292 38966 19348 39004
rect 19180 38770 19236 38780
rect 19068 38724 19124 38734
rect 19404 38668 19460 46732
rect 19964 45892 20020 45902
rect 19964 45798 20020 45836
rect 19628 45556 19684 45566
rect 19628 44548 19684 45500
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19964 44996 20020 45006
rect 20188 44996 20244 49200
rect 19964 44994 20244 44996
rect 19964 44942 19966 44994
rect 20018 44942 20244 44994
rect 19964 44940 20244 44942
rect 20300 47236 20356 47246
rect 20300 46004 20356 47180
rect 19964 44930 20020 44940
rect 19628 44436 19684 44492
rect 19516 44434 19684 44436
rect 19516 44382 19630 44434
rect 19682 44382 19684 44434
rect 19516 44380 19684 44382
rect 19516 42754 19572 44380
rect 19628 44370 19684 44380
rect 20300 44322 20356 45948
rect 20524 47124 20580 47134
rect 20524 44434 20580 47068
rect 21084 46004 21140 46014
rect 20636 45890 20692 45902
rect 20636 45838 20638 45890
rect 20690 45838 20692 45890
rect 20636 45332 20692 45838
rect 20636 45108 20692 45276
rect 20972 45220 21028 45230
rect 20860 45108 20916 45118
rect 20636 45106 20916 45108
rect 20636 45054 20862 45106
rect 20914 45054 20916 45106
rect 20636 45052 20916 45054
rect 20860 44772 20916 45052
rect 20860 44706 20916 44716
rect 20524 44382 20526 44434
rect 20578 44382 20580 44434
rect 20524 44370 20580 44382
rect 20300 44270 20302 44322
rect 20354 44270 20356 44322
rect 20300 44258 20356 44270
rect 20860 44212 20916 44222
rect 20860 44118 20916 44156
rect 20188 44100 20244 44110
rect 20412 44100 20468 44110
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19516 42702 19518 42754
rect 19570 42702 19572 42754
rect 19516 42690 19572 42702
rect 19628 43428 19684 43438
rect 19628 42420 19684 43372
rect 20076 42868 20132 42878
rect 20076 42754 20132 42812
rect 20076 42702 20078 42754
rect 20130 42702 20132 42754
rect 20076 42690 20132 42702
rect 19516 42364 19684 42420
rect 19836 42364 20100 42374
rect 19516 41186 19572 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19964 42084 20020 42094
rect 19516 41134 19518 41186
rect 19570 41134 19572 41186
rect 19516 41122 19572 41134
rect 19852 41858 19908 41870
rect 19852 41806 19854 41858
rect 19906 41806 19908 41858
rect 19852 40964 19908 41806
rect 19964 41186 20020 42028
rect 19964 41134 19966 41186
rect 20018 41134 20020 41186
rect 19964 41122 20020 41134
rect 19852 40898 19908 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19852 40628 19908 40638
rect 19852 40514 19908 40572
rect 19852 40462 19854 40514
rect 19906 40462 19908 40514
rect 19852 40450 19908 40462
rect 20188 40292 20244 44044
rect 20300 44098 20468 44100
rect 20300 44046 20414 44098
rect 20466 44046 20468 44098
rect 20300 44044 20468 44046
rect 20300 41636 20356 44044
rect 20412 44034 20468 44044
rect 20636 44100 20692 44110
rect 20636 44006 20692 44044
rect 20636 43876 20692 43886
rect 20636 43426 20692 43820
rect 20636 43374 20638 43426
rect 20690 43374 20692 43426
rect 20636 43362 20692 43374
rect 20860 42980 20916 42990
rect 20748 42868 20804 42878
rect 20748 42774 20804 42812
rect 20860 42754 20916 42924
rect 20860 42702 20862 42754
rect 20914 42702 20916 42754
rect 20524 42642 20580 42654
rect 20524 42590 20526 42642
rect 20578 42590 20580 42642
rect 20524 42196 20580 42590
rect 20636 42532 20692 42542
rect 20860 42532 20916 42702
rect 20636 42530 20804 42532
rect 20636 42478 20638 42530
rect 20690 42478 20804 42530
rect 20636 42476 20804 42478
rect 20636 42466 20692 42476
rect 20524 42130 20580 42140
rect 20636 42084 20692 42094
rect 20300 41570 20356 41580
rect 20524 41970 20580 41982
rect 20524 41918 20526 41970
rect 20578 41918 20580 41970
rect 20412 41524 20468 41534
rect 19964 40236 20244 40292
rect 20300 41188 20356 41198
rect 20300 40740 20356 41132
rect 19964 39506 20020 40236
rect 20300 40180 20356 40684
rect 20412 41186 20468 41468
rect 20524 41412 20580 41918
rect 20524 41346 20580 41356
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 20412 40404 20468 41134
rect 20524 41188 20580 41198
rect 20636 41188 20692 42028
rect 20748 41860 20804 42476
rect 20860 42466 20916 42476
rect 20972 42084 21028 45164
rect 20748 41794 20804 41804
rect 20860 42028 21028 42084
rect 20860 41524 20916 42028
rect 21084 41972 21140 45948
rect 21308 45890 21364 45902
rect 21308 45838 21310 45890
rect 21362 45838 21364 45890
rect 21308 44772 21364 45838
rect 21420 45108 21476 45118
rect 21420 45014 21476 45052
rect 21308 44706 21364 44716
rect 21196 43428 21252 43438
rect 21196 42980 21252 43372
rect 21532 43428 21588 49200
rect 24220 48244 24276 48254
rect 22092 45890 22148 45902
rect 22092 45838 22094 45890
rect 22146 45838 22148 45890
rect 22092 45556 22148 45838
rect 22092 45490 22148 45500
rect 24220 45444 24276 48188
rect 25452 48132 25508 48142
rect 24892 46564 24948 46574
rect 24444 46452 24500 46462
rect 24444 46002 24500 46396
rect 24444 45950 24446 46002
rect 24498 45950 24500 46002
rect 24444 45938 24500 45950
rect 24668 46116 24724 46126
rect 23772 45332 23828 45342
rect 23772 45238 23828 45276
rect 24220 45106 24276 45388
rect 24444 45556 24500 45566
rect 24444 45330 24500 45500
rect 24444 45278 24446 45330
rect 24498 45278 24500 45330
rect 24444 45266 24500 45278
rect 24556 45108 24612 45118
rect 24220 45054 24222 45106
rect 24274 45054 24276 45106
rect 24220 45042 24276 45054
rect 24332 45106 24612 45108
rect 24332 45054 24558 45106
rect 24610 45054 24612 45106
rect 24332 45052 24612 45054
rect 22316 44660 22372 44670
rect 21644 44322 21700 44334
rect 21644 44270 21646 44322
rect 21698 44270 21700 44322
rect 21644 43540 21700 44270
rect 21644 43474 21700 43484
rect 21980 43540 22036 43550
rect 21532 43362 21588 43372
rect 21196 42914 21252 42924
rect 21644 42868 21700 42878
rect 20860 41458 20916 41468
rect 20972 41916 21140 41972
rect 21308 42866 21700 42868
rect 21308 42814 21646 42866
rect 21698 42814 21700 42866
rect 21308 42812 21700 42814
rect 20524 41186 20636 41188
rect 20524 41134 20526 41186
rect 20578 41134 20636 41186
rect 20524 41132 20636 41134
rect 20524 41122 20580 41132
rect 20636 41122 20692 41132
rect 20748 41076 20804 41086
rect 20636 40964 20692 40974
rect 20748 40964 20804 41020
rect 20636 40962 20804 40964
rect 20636 40910 20638 40962
rect 20690 40910 20804 40962
rect 20636 40908 20804 40910
rect 20636 40898 20692 40908
rect 20972 40628 21028 41916
rect 21196 41860 21252 41870
rect 20412 40338 20468 40348
rect 20636 40572 21028 40628
rect 20636 40402 20692 40572
rect 20636 40350 20638 40402
rect 20690 40350 20692 40402
rect 20636 40338 20692 40350
rect 20748 40404 20804 40414
rect 20188 40124 20356 40180
rect 20188 39618 20244 40124
rect 20300 39732 20356 39742
rect 20300 39638 20356 39676
rect 20188 39566 20190 39618
rect 20242 39566 20244 39618
rect 20188 39554 20244 39566
rect 20412 39620 20468 39630
rect 20636 39620 20692 39630
rect 20412 39618 20636 39620
rect 20412 39566 20414 39618
rect 20466 39566 20636 39618
rect 20412 39564 20636 39566
rect 20412 39554 20468 39564
rect 19964 39454 19966 39506
rect 20018 39454 20020 39506
rect 19964 39396 20020 39454
rect 19964 39340 20244 39396
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 39060 20244 39340
rect 20076 39004 20244 39060
rect 19964 38946 20020 38958
rect 19964 38894 19966 38946
rect 20018 38894 20020 38946
rect 19964 38836 20020 38894
rect 19852 38724 19908 38734
rect 18620 38612 18900 38668
rect 19068 38612 19348 38668
rect 19404 38612 19572 38668
rect 19852 38630 19908 38668
rect 18396 38162 18452 38174
rect 18396 38110 18398 38162
rect 18450 38110 18452 38162
rect 18172 37492 18228 37502
rect 18060 37490 18228 37492
rect 18060 37438 18174 37490
rect 18226 37438 18228 37490
rect 18060 37436 18228 37438
rect 18172 37426 18228 37436
rect 18284 37380 18340 37390
rect 18284 37286 18340 37324
rect 17612 37214 17614 37266
rect 17666 37214 17668 37266
rect 17612 37202 17668 37214
rect 18060 37268 18116 37278
rect 18060 37266 18228 37268
rect 18060 37214 18062 37266
rect 18114 37214 18228 37266
rect 18060 37212 18228 37214
rect 18060 37202 18116 37212
rect 17500 36988 17668 37044
rect 17500 36820 17556 36830
rect 17500 36594 17556 36764
rect 17500 36542 17502 36594
rect 17554 36542 17556 36594
rect 17500 36530 17556 36542
rect 17276 36430 17278 36482
rect 17330 36430 17332 36482
rect 17276 36148 17332 36430
rect 17612 36372 17668 36988
rect 17612 36278 17668 36316
rect 18172 36260 18228 37212
rect 18396 36484 18452 38110
rect 18732 37828 18788 37838
rect 18396 36418 18452 36428
rect 18508 37492 18564 37502
rect 18508 37156 18564 37436
rect 18508 36482 18564 37100
rect 18508 36430 18510 36482
rect 18562 36430 18564 36482
rect 18508 36418 18564 36430
rect 18620 36372 18676 36382
rect 18172 36258 18340 36260
rect 18172 36206 18174 36258
rect 18226 36206 18340 36258
rect 18172 36204 18340 36206
rect 18172 36194 18228 36204
rect 17276 36082 17332 36092
rect 18060 36148 18116 36158
rect 17724 35924 17780 35934
rect 16940 35922 17780 35924
rect 16940 35870 17726 35922
rect 17778 35870 17780 35922
rect 16940 35868 17780 35870
rect 18060 35924 18116 36092
rect 18284 36148 18340 36204
rect 18284 36082 18340 36092
rect 18172 35924 18228 35934
rect 18060 35922 18228 35924
rect 18060 35870 18174 35922
rect 18226 35870 18228 35922
rect 18060 35868 18228 35870
rect 17724 35858 17780 35868
rect 18172 35858 18228 35868
rect 18620 35924 18676 36316
rect 18620 35830 18676 35868
rect 16828 35756 17108 35812
rect 16604 35634 16660 35644
rect 17052 35698 17108 35756
rect 17052 35646 17054 35698
rect 17106 35646 17108 35698
rect 17052 35634 17108 35646
rect 15708 35186 15764 35196
rect 17948 35588 18004 35598
rect 17500 35028 17556 35038
rect 17500 34934 17556 34972
rect 17948 35026 18004 35532
rect 17948 34974 17950 35026
rect 18002 34974 18004 35026
rect 17948 34962 18004 34974
rect 18620 35028 18676 35038
rect 18732 35028 18788 37772
rect 18844 37490 18900 38612
rect 19180 38500 19236 38510
rect 18844 37438 18846 37490
rect 18898 37438 18900 37490
rect 18844 37426 18900 37438
rect 18956 38276 19012 38286
rect 18956 38050 19012 38220
rect 18956 37998 18958 38050
rect 19010 37998 19012 38050
rect 18956 37044 19012 37998
rect 19068 37826 19124 37838
rect 19068 37774 19070 37826
rect 19122 37774 19124 37826
rect 19068 37716 19124 37774
rect 19180 37828 19236 38444
rect 19292 37940 19348 38612
rect 19404 37940 19460 37950
rect 19292 37938 19460 37940
rect 19292 37886 19406 37938
rect 19458 37886 19460 37938
rect 19292 37884 19460 37886
rect 19404 37874 19460 37884
rect 19180 37734 19236 37772
rect 19068 37650 19124 37660
rect 19292 37716 19348 37726
rect 19180 37604 19236 37614
rect 19180 37380 19236 37548
rect 18956 36978 19012 36988
rect 19068 37378 19236 37380
rect 19068 37326 19182 37378
rect 19234 37326 19236 37378
rect 19068 37324 19236 37326
rect 19068 37156 19124 37324
rect 19180 37314 19236 37324
rect 18956 36596 19012 36606
rect 19068 36596 19124 37100
rect 18956 36594 19124 36596
rect 18956 36542 18958 36594
rect 19010 36542 19124 36594
rect 18956 36540 19124 36542
rect 18956 36530 19012 36540
rect 19180 36484 19236 36494
rect 19180 36148 19236 36428
rect 19068 35924 19124 35934
rect 19180 35924 19236 36092
rect 19068 35922 19236 35924
rect 19068 35870 19070 35922
rect 19122 35870 19236 35922
rect 19068 35868 19236 35870
rect 19068 35858 19124 35868
rect 19292 35140 19348 37660
rect 19404 37604 19460 37614
rect 19404 36594 19460 37548
rect 19516 37492 19572 38612
rect 19964 38612 20020 38780
rect 19964 38546 20020 38556
rect 19628 38500 19684 38510
rect 19628 37716 19684 38444
rect 19964 38388 20020 38398
rect 19964 38052 20020 38332
rect 20076 38276 20132 39004
rect 20188 38834 20244 38846
rect 20188 38782 20190 38834
rect 20242 38782 20244 38834
rect 20188 38388 20244 38782
rect 20412 38834 20468 38846
rect 20412 38782 20414 38834
rect 20466 38782 20468 38834
rect 20412 38500 20468 38782
rect 20412 38434 20468 38444
rect 20188 38322 20244 38332
rect 20076 38210 20132 38220
rect 20636 38274 20692 39564
rect 20636 38222 20638 38274
rect 20690 38222 20692 38274
rect 20636 38210 20692 38222
rect 20076 38052 20132 38062
rect 19964 38050 20132 38052
rect 19964 37998 20078 38050
rect 20130 37998 20132 38050
rect 19964 37996 20132 37998
rect 20076 37986 20132 37996
rect 20412 37940 20468 37950
rect 20412 37846 20468 37884
rect 20300 37828 20356 37838
rect 19628 37650 19684 37660
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20300 37604 20356 37772
rect 20300 37548 20468 37604
rect 19852 37492 19908 37502
rect 19516 37490 19908 37492
rect 19516 37438 19854 37490
rect 19906 37438 19908 37490
rect 19516 37436 19908 37438
rect 19852 37426 19908 37436
rect 20076 37492 20132 37502
rect 19740 37156 19796 37166
rect 19740 37062 19796 37100
rect 19404 36542 19406 36594
rect 19458 36542 19460 36594
rect 19404 36530 19460 36542
rect 19516 37044 19572 37054
rect 19516 35922 19572 36988
rect 19964 36260 20020 36336
rect 19516 35870 19518 35922
rect 19570 35870 19572 35922
rect 19516 35474 19572 35870
rect 19516 35422 19518 35474
rect 19570 35422 19572 35474
rect 19516 35410 19572 35422
rect 19628 36204 19964 36260
rect 20076 36260 20132 37436
rect 20300 37156 20356 37166
rect 20300 37062 20356 37100
rect 20412 36594 20468 37548
rect 20524 37380 20580 37390
rect 20524 37044 20580 37324
rect 20524 36978 20580 36988
rect 20412 36542 20414 36594
rect 20466 36542 20468 36594
rect 20412 36530 20468 36542
rect 20076 36204 20244 36260
rect 18620 35026 18788 35028
rect 18620 34974 18622 35026
rect 18674 34974 18788 35026
rect 18620 34972 18788 34974
rect 19068 35084 19348 35140
rect 19068 35026 19124 35084
rect 19068 34974 19070 35026
rect 19122 34974 19124 35026
rect 18620 34962 18676 34972
rect 19068 34962 19124 34974
rect 19628 33572 19684 36204
rect 19964 36194 20020 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19964 35924 20020 35934
rect 20188 35924 20244 36204
rect 19964 35922 20244 35924
rect 19964 35870 19966 35922
rect 20018 35870 20244 35922
rect 19964 35868 20244 35870
rect 20748 35924 20804 40348
rect 20972 40404 21028 40572
rect 20972 40338 21028 40348
rect 21084 41858 21252 41860
rect 21084 41806 21198 41858
rect 21250 41806 21252 41858
rect 21084 41804 21252 41806
rect 20860 40068 20916 40078
rect 20860 39732 20916 40012
rect 20860 39730 21028 39732
rect 20860 39678 20862 39730
rect 20914 39678 21028 39730
rect 20860 39676 21028 39678
rect 20860 39666 20916 39676
rect 20972 38946 21028 39676
rect 20972 38894 20974 38946
rect 21026 38894 21028 38946
rect 20972 38882 21028 38894
rect 20860 38724 20916 38734
rect 20860 38612 21028 38668
rect 20860 38388 20916 38398
rect 20860 37826 20916 38332
rect 20860 37774 20862 37826
rect 20914 37774 20916 37826
rect 20860 37380 20916 37774
rect 20972 37492 21028 38612
rect 21084 38500 21140 41804
rect 21196 41794 21252 41804
rect 21196 41188 21252 41198
rect 21196 40514 21252 41132
rect 21196 40462 21198 40514
rect 21250 40462 21252 40514
rect 21196 40450 21252 40462
rect 21308 40180 21364 42812
rect 21644 42802 21700 42812
rect 21756 42196 21812 42206
rect 21644 41188 21700 41198
rect 21532 41186 21700 41188
rect 21532 41134 21646 41186
rect 21698 41134 21700 41186
rect 21532 41132 21700 41134
rect 21084 38434 21140 38444
rect 21196 40124 21364 40180
rect 21420 40402 21476 40414
rect 21420 40350 21422 40402
rect 21474 40350 21476 40402
rect 21084 38274 21140 38286
rect 21084 38222 21086 38274
rect 21138 38222 21140 38274
rect 21084 37492 21140 38222
rect 21196 37716 21252 40124
rect 21308 39844 21364 39854
rect 21308 39058 21364 39788
rect 21308 39006 21310 39058
rect 21362 39006 21364 39058
rect 21308 38724 21364 39006
rect 21420 38836 21476 40350
rect 21532 38948 21588 41132
rect 21644 41122 21700 41132
rect 21756 41186 21812 42140
rect 21756 41134 21758 41186
rect 21810 41134 21812 41186
rect 21756 41122 21812 41134
rect 21868 40962 21924 40974
rect 21868 40910 21870 40962
rect 21922 40910 21924 40962
rect 21644 40852 21700 40862
rect 21644 40626 21700 40796
rect 21644 40574 21646 40626
rect 21698 40574 21700 40626
rect 21644 40562 21700 40574
rect 21756 40402 21812 40414
rect 21756 40350 21758 40402
rect 21810 40350 21812 40402
rect 21756 40180 21812 40350
rect 21756 40114 21812 40124
rect 21868 39844 21924 40910
rect 21868 39778 21924 39788
rect 21980 39732 22036 43484
rect 22092 41860 22148 41870
rect 22092 41076 22148 41804
rect 22092 41010 22148 41020
rect 22316 40740 22372 44604
rect 22428 44436 22484 44446
rect 22428 44210 22484 44380
rect 22428 44158 22430 44210
rect 22482 44158 22484 44210
rect 22428 43988 22484 44158
rect 22428 43922 22484 43932
rect 24108 43540 24164 43550
rect 24332 43540 24388 45052
rect 24556 45042 24612 45052
rect 24444 44548 24500 44558
rect 24444 43652 24500 44492
rect 24556 44436 24612 44446
rect 24668 44436 24724 46060
rect 24556 44434 24668 44436
rect 24556 44382 24558 44434
rect 24610 44382 24668 44434
rect 24556 44380 24668 44382
rect 24556 44370 24612 44380
rect 24668 44304 24724 44380
rect 24780 45106 24836 45118
rect 24780 45054 24782 45106
rect 24834 45054 24836 45106
rect 24444 43586 24500 43596
rect 24556 44100 24612 44110
rect 24556 43650 24612 44044
rect 24780 43876 24836 45054
rect 24556 43598 24558 43650
rect 24610 43598 24612 43650
rect 24556 43586 24612 43598
rect 24668 43820 24836 43876
rect 24108 43538 24388 43540
rect 24108 43486 24110 43538
rect 24162 43486 24388 43538
rect 24108 43484 24388 43486
rect 24108 43474 24164 43484
rect 22316 40626 22372 40684
rect 22316 40574 22318 40626
rect 22370 40574 22372 40626
rect 22316 40404 22372 40574
rect 22316 40338 22372 40348
rect 22428 43428 22484 43438
rect 23324 43428 23380 43438
rect 22204 40178 22260 40190
rect 22204 40126 22206 40178
rect 22258 40126 22260 40178
rect 22204 40068 22260 40126
rect 22204 40002 22260 40012
rect 21980 39676 22148 39732
rect 21644 39508 21700 39518
rect 21644 39414 21700 39452
rect 21980 39508 22036 39518
rect 21980 39414 22036 39452
rect 21868 39172 21924 39182
rect 21868 39058 21924 39116
rect 21868 39006 21870 39058
rect 21922 39006 21924 39058
rect 21532 38892 21812 38948
rect 21420 38770 21476 38780
rect 21308 38658 21364 38668
rect 21532 38724 21588 38734
rect 21532 38612 21700 38668
rect 21532 38388 21588 38398
rect 21532 38162 21588 38332
rect 21532 38110 21534 38162
rect 21586 38110 21588 38162
rect 21532 38098 21588 38110
rect 21196 37660 21476 37716
rect 21196 37492 21252 37502
rect 21084 37490 21252 37492
rect 21084 37438 21198 37490
rect 21250 37438 21252 37490
rect 21084 37436 21252 37438
rect 20972 37426 21028 37436
rect 20860 37314 20916 37324
rect 20860 37154 20916 37166
rect 20860 37102 20862 37154
rect 20914 37102 20916 37154
rect 20860 37044 20916 37102
rect 20860 36978 20916 36988
rect 20972 37156 21028 37166
rect 20972 36594 21028 37100
rect 20972 36542 20974 36594
rect 21026 36542 21028 36594
rect 20972 36530 21028 36542
rect 20860 35924 20916 35934
rect 20748 35922 20916 35924
rect 20748 35870 20862 35922
rect 20914 35870 20916 35922
rect 20748 35868 20916 35870
rect 19964 35858 20020 35868
rect 20860 35858 20916 35868
rect 21196 35700 21252 37436
rect 21420 36596 21476 37660
rect 21644 37492 21700 38612
rect 21756 37828 21812 38892
rect 21756 37762 21812 37772
rect 21756 37492 21812 37502
rect 21644 37490 21812 37492
rect 21644 37438 21758 37490
rect 21810 37438 21812 37490
rect 21644 37436 21812 37438
rect 21756 37426 21812 37436
rect 21532 36596 21588 36606
rect 21420 36594 21588 36596
rect 21420 36542 21534 36594
rect 21586 36542 21588 36594
rect 21420 36540 21588 36542
rect 21420 35924 21476 36540
rect 21532 36530 21588 36540
rect 21420 35858 21476 35868
rect 21196 35634 21252 35644
rect 20412 35586 20468 35598
rect 20412 35534 20414 35586
rect 20466 35534 20468 35586
rect 20412 35474 20468 35534
rect 20412 35422 20414 35474
rect 20466 35422 20468 35474
rect 20412 35410 20468 35422
rect 21868 35028 21924 39006
rect 21980 38948 22036 38958
rect 22092 38948 22148 39676
rect 21980 38946 22148 38948
rect 21980 38894 21982 38946
rect 22034 38894 22094 38946
rect 22146 38894 22148 38946
rect 21980 38892 22148 38894
rect 21980 38882 22036 38892
rect 22092 38816 22148 38892
rect 22204 39508 22260 39518
rect 22428 39508 22484 43372
rect 23212 43426 23380 43428
rect 23212 43374 23326 43426
rect 23378 43374 23380 43426
rect 23212 43372 23380 43374
rect 22876 43204 22932 43214
rect 22764 41524 22820 41534
rect 22764 41074 22820 41468
rect 22764 41022 22766 41074
rect 22818 41022 22820 41074
rect 22764 41010 22820 41022
rect 22652 40962 22708 40974
rect 22652 40910 22654 40962
rect 22706 40910 22708 40962
rect 22540 40516 22596 40526
rect 22540 40422 22596 40460
rect 22540 39508 22596 39518
rect 22428 39506 22596 39508
rect 22428 39454 22542 39506
rect 22594 39454 22596 39506
rect 22428 39452 22596 39454
rect 22092 38164 22148 38174
rect 22204 38164 22260 39452
rect 22540 39442 22596 39452
rect 22428 39058 22484 39070
rect 22428 39006 22430 39058
rect 22482 39006 22484 39058
rect 22092 38162 22260 38164
rect 22092 38110 22094 38162
rect 22146 38110 22260 38162
rect 22092 38108 22260 38110
rect 22316 38948 22372 38958
rect 22428 38948 22484 39006
rect 22652 39060 22708 40910
rect 22652 38994 22708 39004
rect 22764 40404 22820 40414
rect 22764 39618 22820 40348
rect 22764 39566 22766 39618
rect 22818 39566 22820 39618
rect 22316 38946 22484 38948
rect 22316 38894 22318 38946
rect 22370 38894 22484 38946
rect 22316 38892 22484 38894
rect 22092 38098 22148 38108
rect 22092 37828 22148 37838
rect 22092 37490 22148 37772
rect 22092 37438 22094 37490
rect 22146 37438 22148 37490
rect 22092 36932 22148 37438
rect 22092 36866 22148 36876
rect 22092 36596 22148 36606
rect 22316 36596 22372 38892
rect 22764 38724 22820 39566
rect 22764 38658 22820 38668
rect 22876 40402 22932 43148
rect 23212 41636 23268 43372
rect 23324 43362 23380 43372
rect 24220 43316 24276 43326
rect 24108 43092 24164 43102
rect 23436 42980 23492 42990
rect 23212 41570 23268 41580
rect 23324 41858 23380 41870
rect 23324 41806 23326 41858
rect 23378 41806 23380 41858
rect 23212 41188 23268 41198
rect 23212 41094 23268 41132
rect 22988 40962 23044 40974
rect 22988 40910 22990 40962
rect 23042 40910 23044 40962
rect 22988 40740 23044 40910
rect 22988 40674 23044 40684
rect 22876 40350 22878 40402
rect 22930 40350 22932 40402
rect 22428 38276 22484 38286
rect 22428 38162 22484 38220
rect 22876 38276 22932 40350
rect 23100 40516 23156 40526
rect 23324 40516 23380 41806
rect 23100 39842 23156 40460
rect 23100 39790 23102 39842
rect 23154 39790 23156 39842
rect 23100 39778 23156 39790
rect 23212 40460 23380 40516
rect 22988 39618 23044 39630
rect 22988 39566 22990 39618
rect 23042 39566 23044 39618
rect 22988 39508 23044 39566
rect 23100 39508 23156 39518
rect 22988 39506 23156 39508
rect 22988 39454 23102 39506
rect 23154 39454 23156 39506
rect 22988 39452 23156 39454
rect 23100 39442 23156 39452
rect 22988 38836 23044 38846
rect 22988 38742 23044 38780
rect 22876 38210 22932 38220
rect 22428 38110 22430 38162
rect 22482 38110 22484 38162
rect 22428 38098 22484 38110
rect 22764 38164 22820 38174
rect 22092 36594 22372 36596
rect 22092 36542 22094 36594
rect 22146 36542 22372 36594
rect 22092 36540 22372 36542
rect 22540 37492 22596 37502
rect 22764 37492 22820 38108
rect 22988 38164 23044 38174
rect 22988 38070 23044 38108
rect 23212 37940 23268 40460
rect 23436 40404 23492 42924
rect 23772 42644 23828 42654
rect 23660 42642 23828 42644
rect 23660 42590 23774 42642
rect 23826 42590 23828 42642
rect 23660 42588 23828 42590
rect 23324 40348 23492 40404
rect 23548 41636 23604 41646
rect 23548 40404 23604 41580
rect 23324 40290 23380 40348
rect 23324 40238 23326 40290
rect 23378 40238 23380 40290
rect 23324 40226 23380 40238
rect 23436 40180 23492 40190
rect 23548 40180 23604 40348
rect 23436 40178 23604 40180
rect 23436 40126 23438 40178
rect 23490 40126 23604 40178
rect 23436 40124 23604 40126
rect 23436 40114 23492 40124
rect 23324 39842 23380 39854
rect 23324 39790 23326 39842
rect 23378 39790 23380 39842
rect 23324 39058 23380 39790
rect 23548 39842 23604 39854
rect 23548 39790 23550 39842
rect 23602 39790 23604 39842
rect 23548 39730 23604 39790
rect 23548 39678 23550 39730
rect 23602 39678 23604 39730
rect 23548 39666 23604 39678
rect 23324 39006 23326 39058
rect 23378 39006 23380 39058
rect 23324 38994 23380 39006
rect 23660 38668 23716 42588
rect 23772 42578 23828 42588
rect 24108 42420 24164 43036
rect 24108 42354 24164 42364
rect 24108 41970 24164 41982
rect 24108 41918 24110 41970
rect 24162 41918 24164 41970
rect 23996 41524 24052 41534
rect 23996 41188 24052 41468
rect 23884 41186 24052 41188
rect 23884 41134 23998 41186
rect 24050 41134 24052 41186
rect 23884 41132 24052 41134
rect 23772 41076 23828 41086
rect 23772 40982 23828 41020
rect 23772 40180 23828 40190
rect 23772 39058 23828 40124
rect 23884 39842 23940 41132
rect 23996 41122 24052 41132
rect 24108 41076 24164 41918
rect 23996 40964 24052 40974
rect 23996 40626 24052 40908
rect 24108 40852 24164 41020
rect 24108 40786 24164 40796
rect 23996 40574 23998 40626
rect 24050 40574 24052 40626
rect 23996 40562 24052 40574
rect 24220 40628 24276 43260
rect 24332 40852 24388 43484
rect 24556 42756 24612 42766
rect 24556 42662 24612 42700
rect 24668 42084 24724 43820
rect 24780 43652 24836 43662
rect 24780 42308 24836 43596
rect 24892 43650 24948 46508
rect 25340 46004 25396 46014
rect 25340 45910 25396 45948
rect 25228 45892 25284 45902
rect 24892 43598 24894 43650
rect 24946 43598 24948 43650
rect 24892 42980 24948 43598
rect 24892 42914 24948 42924
rect 25004 44436 25060 44446
rect 25004 43316 25060 44380
rect 25228 44434 25284 45836
rect 25228 44382 25230 44434
rect 25282 44382 25284 44434
rect 25228 44370 25284 44382
rect 25340 44772 25396 44782
rect 25116 44098 25172 44110
rect 25340 44100 25396 44716
rect 25116 44046 25118 44098
rect 25170 44046 25172 44098
rect 25116 43764 25172 44046
rect 25116 43698 25172 43708
rect 25228 44098 25396 44100
rect 25228 44046 25342 44098
rect 25394 44046 25396 44098
rect 25228 44044 25396 44046
rect 25004 42756 25060 43260
rect 25004 42690 25060 42700
rect 25116 43092 25172 43102
rect 25116 42642 25172 43036
rect 25116 42590 25118 42642
rect 25170 42590 25172 42642
rect 25116 42578 25172 42590
rect 25004 42532 25060 42542
rect 25004 42438 25060 42476
rect 24780 42252 25172 42308
rect 24668 42028 24948 42084
rect 24780 41860 24836 41870
rect 24780 41766 24836 41804
rect 24668 41746 24724 41758
rect 24668 41694 24670 41746
rect 24722 41694 24724 41746
rect 24668 41524 24724 41694
rect 24668 41458 24724 41468
rect 24780 41412 24836 41422
rect 24780 41298 24836 41356
rect 24780 41246 24782 41298
rect 24834 41246 24836 41298
rect 24780 41234 24836 41246
rect 24892 41076 24948 42028
rect 24780 41020 24948 41076
rect 25004 41524 25060 41534
rect 24332 40786 24388 40796
rect 24668 40962 24724 40974
rect 24668 40910 24670 40962
rect 24722 40910 24724 40962
rect 24668 40740 24724 40910
rect 24668 40674 24724 40684
rect 24556 40628 24612 40638
rect 24220 40626 24612 40628
rect 24220 40574 24558 40626
rect 24610 40574 24612 40626
rect 24220 40572 24612 40574
rect 24108 40516 24164 40526
rect 24220 40516 24276 40572
rect 24556 40562 24612 40572
rect 24108 40514 24276 40516
rect 24108 40462 24110 40514
rect 24162 40462 24276 40514
rect 24108 40460 24276 40462
rect 24108 40450 24164 40460
rect 23996 40404 24052 40414
rect 24780 40404 24836 41020
rect 23996 40292 24052 40348
rect 24668 40348 24836 40404
rect 23996 40236 24276 40292
rect 23884 39790 23886 39842
rect 23938 39790 23940 39842
rect 23884 39778 23940 39790
rect 23996 39620 24052 39630
rect 23996 39526 24052 39564
rect 23772 39006 23774 39058
rect 23826 39006 23828 39058
rect 23772 38994 23828 39006
rect 23436 38612 23716 38668
rect 23436 38052 23492 38612
rect 24220 38164 24276 40236
rect 24444 39842 24500 39854
rect 24444 39790 24446 39842
rect 24498 39790 24500 39842
rect 24444 39730 24500 39790
rect 24444 39678 24446 39730
rect 24498 39678 24500 39730
rect 24444 39666 24500 39678
rect 24332 39396 24388 39406
rect 24332 39060 24388 39340
rect 24332 38966 24388 39004
rect 24668 39058 24724 40348
rect 25004 40292 25060 41468
rect 24668 39006 24670 39058
rect 24722 39006 24724 39058
rect 24332 38164 24388 38174
rect 24220 38162 24388 38164
rect 24220 38110 24334 38162
rect 24386 38110 24388 38162
rect 24220 38108 24388 38110
rect 24332 38098 24388 38108
rect 23436 37958 23492 37996
rect 23212 37874 23268 37884
rect 23772 37826 23828 37838
rect 23772 37774 23774 37826
rect 23826 37774 23828 37826
rect 22988 37492 23044 37502
rect 22764 37436 22988 37492
rect 22092 36530 22148 36540
rect 22540 35588 22596 37436
rect 22988 37398 23044 37436
rect 23772 36820 23828 37774
rect 23772 36754 23828 36764
rect 24668 36372 24724 39006
rect 24780 40236 25060 40292
rect 24780 37716 24836 40236
rect 24780 37650 24836 37660
rect 24892 40068 24948 40078
rect 24892 37492 24948 40012
rect 25004 39732 25060 39742
rect 25116 39732 25172 42252
rect 25004 39730 25172 39732
rect 25004 39678 25006 39730
rect 25058 39678 25172 39730
rect 25004 39676 25172 39678
rect 25004 39666 25060 39676
rect 25116 39620 25172 39676
rect 25116 39554 25172 39564
rect 25228 41524 25284 44044
rect 25340 44034 25396 44044
rect 25452 43092 25508 48076
rect 25676 46340 25732 46350
rect 25452 43026 25508 43036
rect 25564 45106 25620 45118
rect 25564 45054 25566 45106
rect 25618 45054 25620 45106
rect 25564 44098 25620 45054
rect 25564 44046 25566 44098
rect 25618 44046 25620 44098
rect 25564 42868 25620 44046
rect 25676 43764 25732 46284
rect 25900 45780 25956 45790
rect 25788 43764 25844 43774
rect 25676 43762 25844 43764
rect 25676 43710 25790 43762
rect 25842 43710 25844 43762
rect 25676 43708 25844 43710
rect 25788 43698 25844 43708
rect 25564 42802 25620 42812
rect 25676 43538 25732 43550
rect 25676 43486 25678 43538
rect 25730 43486 25732 43538
rect 25564 42644 25620 42682
rect 25564 42578 25620 42588
rect 25340 42532 25396 42542
rect 25452 42532 25508 42542
rect 25340 42530 25452 42532
rect 25340 42478 25342 42530
rect 25394 42478 25452 42530
rect 25340 42476 25452 42478
rect 25340 42466 25396 42476
rect 24892 37426 24948 37436
rect 25228 36484 25284 41468
rect 25340 41860 25396 41870
rect 25340 41298 25396 41804
rect 25340 41246 25342 41298
rect 25394 41246 25396 41298
rect 25340 41234 25396 41246
rect 25340 40852 25396 40862
rect 25340 40068 25396 40796
rect 25340 40002 25396 40012
rect 25452 40852 25508 42476
rect 25564 42420 25620 42430
rect 25564 41410 25620 42364
rect 25676 42084 25732 43486
rect 25676 42018 25732 42028
rect 25788 41972 25844 41982
rect 25900 41972 25956 45724
rect 26908 45780 26964 49200
rect 29372 48020 29428 48030
rect 26908 45714 26964 45724
rect 27020 47908 27076 47918
rect 26236 45668 26292 45678
rect 26236 45330 26292 45612
rect 26236 45278 26238 45330
rect 26290 45278 26292 45330
rect 26236 45266 26292 45278
rect 27020 45330 27076 47852
rect 27356 47572 27412 47582
rect 27244 47348 27300 47358
rect 27020 45278 27022 45330
rect 27074 45278 27076 45330
rect 27020 45266 27076 45278
rect 27132 46228 27188 46238
rect 27132 45556 27188 46172
rect 27132 45218 27188 45500
rect 27132 45166 27134 45218
rect 27186 45166 27188 45218
rect 27132 45154 27188 45166
rect 26012 45106 26068 45118
rect 26012 45054 26014 45106
rect 26066 45054 26068 45106
rect 26012 44772 26068 45054
rect 26124 45108 26180 45118
rect 26684 45108 26740 45118
rect 26124 45014 26180 45052
rect 26572 45106 26740 45108
rect 26572 45054 26686 45106
rect 26738 45054 26740 45106
rect 26572 45052 26740 45054
rect 26572 44996 26628 45052
rect 26684 45042 26740 45052
rect 26012 44706 26068 44716
rect 26348 44940 26628 44996
rect 26236 44212 26292 44222
rect 26236 44118 26292 44156
rect 26012 44100 26068 44110
rect 26012 43650 26068 44044
rect 26012 43598 26014 43650
rect 26066 43598 26068 43650
rect 26012 43586 26068 43598
rect 26236 43538 26292 43550
rect 26236 43486 26238 43538
rect 26290 43486 26292 43538
rect 25788 41970 25956 41972
rect 25788 41918 25790 41970
rect 25842 41918 25902 41970
rect 25954 41918 25956 41970
rect 25788 41916 25956 41918
rect 25788 41906 25844 41916
rect 25900 41840 25956 41916
rect 26012 43316 26068 43326
rect 25564 41358 25566 41410
rect 25618 41358 25620 41410
rect 25564 41346 25620 41358
rect 25676 41746 25732 41758
rect 25676 41694 25678 41746
rect 25730 41694 25732 41746
rect 25676 41300 25732 41694
rect 25676 41234 25732 41244
rect 25788 40962 25844 40974
rect 25788 40910 25790 40962
rect 25842 40910 25844 40962
rect 25788 40852 25844 40910
rect 25452 40796 25844 40852
rect 25340 39844 25396 39854
rect 25340 39730 25396 39788
rect 25340 39678 25342 39730
rect 25394 39678 25396 39730
rect 25340 39666 25396 39678
rect 25452 39508 25508 40796
rect 26012 40740 26068 43260
rect 26236 42756 26292 43486
rect 26348 43428 26404 44940
rect 26684 44884 26740 44894
rect 26572 44212 26628 44222
rect 26684 44212 26740 44828
rect 26796 44324 26852 44334
rect 27244 44324 27300 47292
rect 27356 45220 27412 47516
rect 29036 47460 29092 47470
rect 28364 47236 28420 47246
rect 27468 46788 27524 46798
rect 27468 46116 27524 46732
rect 27468 46002 27524 46060
rect 27468 45950 27470 46002
rect 27522 45950 27524 46002
rect 27468 45938 27524 45950
rect 28252 46564 28308 46574
rect 28252 45892 28308 46508
rect 28252 45798 28308 45836
rect 27356 45126 27412 45164
rect 27916 45106 27972 45118
rect 27916 45054 27918 45106
rect 27970 45054 27972 45106
rect 27692 44884 27748 44894
rect 27692 44436 27748 44828
rect 27356 44324 27412 44334
rect 27244 44268 27356 44324
rect 26796 44230 26852 44268
rect 26572 44210 26740 44212
rect 26572 44158 26574 44210
rect 26626 44158 26740 44210
rect 27356 44192 27412 44268
rect 27692 44210 27748 44380
rect 26572 44156 26740 44158
rect 26572 44146 26628 44156
rect 26348 43362 26404 43372
rect 26460 44098 26516 44110
rect 26460 44046 26462 44098
rect 26514 44046 26516 44098
rect 26460 42868 26516 44046
rect 26684 44100 26740 44156
rect 27692 44158 27694 44210
rect 27746 44158 27748 44210
rect 27692 44146 27748 44158
rect 26460 42812 26628 42868
rect 26124 42532 26180 42542
rect 26124 42438 26180 42476
rect 26236 42084 26292 42700
rect 26460 42642 26516 42654
rect 26460 42590 26462 42642
rect 26514 42590 26516 42642
rect 26236 42028 26404 42084
rect 26124 41972 26180 41982
rect 26124 41970 26292 41972
rect 26124 41918 26126 41970
rect 26178 41918 26292 41970
rect 26124 41916 26292 41918
rect 26124 41906 26180 41916
rect 26236 41858 26292 41916
rect 26236 41806 26238 41858
rect 26290 41806 26292 41858
rect 26236 41794 26292 41806
rect 26236 41188 26292 41198
rect 26236 41094 26292 41132
rect 25564 40684 26068 40740
rect 25564 40626 25620 40684
rect 25564 40574 25566 40626
rect 25618 40574 25620 40626
rect 25564 40562 25620 40574
rect 26012 40404 26068 40414
rect 26012 40310 26068 40348
rect 26348 40180 26404 42028
rect 26460 41748 26516 42590
rect 26460 41682 26516 41692
rect 26460 40852 26516 40862
rect 26460 40626 26516 40796
rect 26460 40574 26462 40626
rect 26514 40574 26516 40626
rect 26460 40562 26516 40574
rect 26348 40114 26404 40124
rect 25788 39620 25844 39630
rect 25788 39526 25844 39564
rect 25452 39442 25508 39452
rect 25228 36418 25284 36428
rect 26236 39394 26292 39406
rect 26236 39342 26238 39394
rect 26290 39342 26292 39394
rect 24668 36306 24724 36316
rect 22540 35522 22596 35532
rect 26236 35252 26292 39342
rect 26572 37044 26628 42812
rect 26684 42644 26740 44044
rect 27692 43764 27748 43774
rect 26796 43540 26852 43550
rect 26908 43540 26964 43550
rect 26852 43538 26964 43540
rect 26852 43486 26910 43538
rect 26962 43486 26964 43538
rect 26852 43484 26964 43486
rect 26796 43474 26852 43484
rect 26908 43474 26964 43484
rect 27132 43540 27188 43550
rect 27244 43540 27300 43550
rect 27132 43538 27244 43540
rect 27132 43486 27134 43538
rect 27186 43486 27244 43538
rect 27132 43484 27244 43486
rect 27132 43474 27188 43484
rect 26684 42578 26740 42588
rect 26796 43314 26852 43326
rect 26796 43262 26798 43314
rect 26850 43262 26852 43314
rect 26796 42532 26852 43262
rect 27020 42980 27076 42990
rect 27020 42886 27076 42924
rect 27132 42868 27188 42878
rect 26684 41858 26740 41870
rect 26684 41806 26686 41858
rect 26738 41806 26740 41858
rect 26684 41748 26740 41806
rect 26684 41682 26740 41692
rect 26684 41410 26740 41422
rect 26684 41358 26686 41410
rect 26738 41358 26740 41410
rect 26684 41298 26740 41358
rect 26684 41246 26686 41298
rect 26738 41246 26740 41298
rect 26684 41234 26740 41246
rect 26572 36978 26628 36988
rect 26796 35812 26852 42476
rect 27020 42644 27076 42654
rect 26908 42420 26964 42430
rect 26908 40626 26964 42364
rect 26908 40574 26910 40626
rect 26962 40574 26964 40626
rect 26908 40562 26964 40574
rect 27020 41860 27076 42588
rect 27132 42196 27188 42812
rect 27244 42644 27300 43484
rect 27692 43426 27748 43708
rect 27916 43652 27972 45054
rect 28140 45106 28196 45118
rect 28140 45054 28142 45106
rect 28194 45054 28196 45106
rect 27804 43540 27860 43550
rect 27804 43446 27860 43484
rect 27692 43374 27694 43426
rect 27746 43374 27748 43426
rect 27580 42868 27636 42878
rect 27580 42774 27636 42812
rect 27468 42756 27524 42766
rect 27244 42588 27412 42644
rect 27132 42140 27300 42196
rect 27132 41860 27188 41870
rect 27020 41858 27188 41860
rect 27020 41806 27134 41858
rect 27186 41806 27188 41858
rect 27020 41804 27188 41806
rect 27020 41746 27076 41804
rect 27132 41794 27188 41804
rect 27020 41694 27022 41746
rect 27074 41694 27076 41746
rect 27020 38836 27076 41694
rect 27244 41298 27300 42140
rect 27244 41246 27246 41298
rect 27298 41246 27300 41298
rect 27244 41234 27300 41246
rect 27356 41076 27412 42588
rect 27020 38770 27076 38780
rect 27132 41020 27412 41076
rect 27132 38668 27188 41020
rect 27356 40628 27412 40638
rect 27356 40534 27412 40572
rect 27020 38612 27188 38668
rect 27020 38388 27076 38612
rect 27020 38322 27076 38332
rect 27468 36596 27524 42700
rect 27692 42644 27748 43374
rect 27916 43204 27972 43596
rect 27916 43138 27972 43148
rect 28028 44994 28084 45006
rect 28028 44942 28030 44994
rect 28082 44942 28084 44994
rect 28028 42868 28084 44942
rect 28140 44660 28196 45054
rect 28364 44996 28420 47180
rect 28364 44930 28420 44940
rect 28476 45106 28532 45118
rect 28476 45054 28478 45106
rect 28530 45054 28532 45106
rect 28140 44100 28196 44604
rect 28364 44660 28420 44670
rect 28364 44322 28420 44604
rect 28364 44270 28366 44322
rect 28418 44270 28420 44322
rect 28364 44258 28420 44270
rect 28140 44034 28196 44044
rect 28028 42802 28084 42812
rect 28140 43876 28196 43886
rect 27580 42588 27748 42644
rect 27580 42420 27636 42588
rect 28028 42532 28084 42542
rect 28028 42438 28084 42476
rect 27580 42364 27972 42420
rect 27692 42196 27748 42206
rect 27580 41858 27636 41870
rect 27580 41806 27582 41858
rect 27634 41806 27636 41858
rect 27580 41746 27636 41806
rect 27580 41694 27582 41746
rect 27634 41694 27636 41746
rect 27580 41682 27636 41694
rect 27692 41298 27748 42140
rect 27692 41246 27694 41298
rect 27746 41246 27748 41298
rect 27692 41234 27748 41246
rect 27916 36820 27972 42364
rect 28028 41858 28084 41870
rect 28028 41806 28030 41858
rect 28082 41806 28084 41858
rect 28028 41524 28084 41806
rect 28028 41458 28084 41468
rect 28028 41300 28084 41310
rect 28140 41300 28196 43820
rect 28476 43764 28532 45054
rect 29036 44994 29092 47404
rect 29260 45778 29316 45790
rect 29260 45726 29262 45778
rect 29314 45726 29316 45778
rect 29036 44942 29038 44994
rect 29090 44942 29092 44994
rect 29036 44930 29092 44942
rect 29148 45218 29204 45230
rect 29148 45166 29150 45218
rect 29202 45166 29204 45218
rect 28924 44660 28980 44670
rect 28588 44100 28644 44110
rect 28588 44006 28644 44044
rect 28252 43708 28532 43764
rect 28588 43876 28644 43886
rect 28252 42308 28308 43708
rect 28476 43540 28532 43550
rect 28588 43540 28644 43820
rect 28924 43764 28980 44604
rect 28924 43650 28980 43708
rect 28924 43598 28926 43650
rect 28978 43598 28980 43650
rect 28924 43586 28980 43598
rect 29148 43876 29204 45166
rect 29260 44548 29316 45726
rect 29372 45218 29428 47964
rect 30044 47796 30100 47806
rect 29372 45166 29374 45218
rect 29426 45166 29428 45218
rect 29372 45108 29428 45166
rect 29372 45042 29428 45052
rect 29484 45778 29540 45790
rect 29484 45726 29486 45778
rect 29538 45726 29540 45778
rect 29372 44548 29428 44558
rect 29260 44492 29372 44548
rect 29372 44212 29428 44492
rect 29484 44436 29540 45726
rect 29820 45778 29876 45790
rect 29820 45726 29822 45778
rect 29874 45726 29876 45778
rect 29596 45668 29652 45678
rect 29596 45574 29652 45612
rect 29484 44370 29540 44380
rect 29596 44996 29652 45006
rect 29484 44212 29540 44222
rect 29372 44210 29540 44212
rect 29372 44158 29486 44210
rect 29538 44158 29540 44210
rect 29372 44156 29540 44158
rect 28476 43538 28644 43540
rect 28476 43486 28478 43538
rect 28530 43486 28644 43538
rect 28476 43484 28644 43486
rect 28476 43474 28532 43484
rect 28364 43426 28420 43438
rect 28364 43374 28366 43426
rect 28418 43374 28420 43426
rect 28364 43316 28420 43374
rect 28364 43250 28420 43260
rect 29148 43204 29204 43820
rect 29372 43540 29428 43550
rect 29372 43446 29428 43484
rect 28924 43148 29148 43204
rect 28476 43092 28532 43102
rect 28476 42866 28532 43036
rect 28476 42814 28478 42866
rect 28530 42814 28532 42866
rect 28476 42802 28532 42814
rect 28252 42242 28308 42252
rect 28924 41970 28980 43148
rect 29148 43138 29204 43148
rect 29484 42868 29540 44156
rect 28924 41918 28926 41970
rect 28978 41918 28980 41970
rect 28924 41906 28980 41918
rect 29372 42812 29540 42868
rect 29372 41970 29428 42812
rect 29484 42530 29540 42542
rect 29484 42478 29486 42530
rect 29538 42478 29540 42530
rect 29484 42308 29540 42478
rect 29484 42242 29540 42252
rect 29596 42196 29652 44940
rect 29820 44212 29876 45726
rect 30044 45220 30100 47740
rect 30940 46228 30996 49200
rect 30940 46172 31444 46228
rect 31388 45890 31444 46172
rect 32284 46004 32340 49200
rect 33180 47124 33236 47134
rect 32284 45938 32340 45948
rect 32396 46116 32452 46126
rect 32396 46002 32452 46060
rect 32396 45950 32398 46002
rect 32450 45950 32452 46002
rect 32396 45938 32452 45950
rect 31388 45838 31390 45890
rect 31442 45838 31444 45890
rect 30380 45780 30436 45790
rect 31164 45780 31220 45790
rect 30380 45686 30436 45724
rect 30940 45778 31220 45780
rect 30940 45726 31166 45778
rect 31218 45726 31220 45778
rect 30940 45724 31220 45726
rect 30604 45556 30660 45566
rect 30044 45218 30212 45220
rect 30044 45166 30046 45218
rect 30098 45166 30212 45218
rect 30044 45164 30212 45166
rect 30044 45154 30100 45164
rect 29932 44996 29988 45006
rect 29932 44902 29988 44940
rect 29932 44324 29988 44334
rect 29932 44230 29988 44268
rect 29820 44146 29876 44156
rect 30044 44212 30100 44222
rect 29820 43426 29876 43438
rect 29820 43374 29822 43426
rect 29874 43374 29876 43426
rect 29820 43316 29876 43374
rect 29820 43250 29876 43260
rect 29932 42868 29988 42878
rect 30044 42868 30100 44156
rect 29932 42866 30100 42868
rect 29932 42814 29934 42866
rect 29986 42814 30100 42866
rect 29932 42812 30100 42814
rect 30156 42868 30212 45164
rect 30604 45218 30660 45500
rect 30716 45444 30772 45454
rect 30716 45330 30772 45388
rect 30716 45278 30718 45330
rect 30770 45278 30772 45330
rect 30716 45266 30772 45278
rect 30604 45166 30606 45218
rect 30658 45166 30660 45218
rect 30604 45154 30660 45166
rect 30828 44660 30884 44670
rect 30828 44434 30884 44604
rect 30828 44382 30830 44434
rect 30882 44382 30884 44434
rect 30828 44370 30884 44382
rect 30380 44212 30436 44222
rect 30380 44118 30436 44156
rect 30716 44100 30772 44110
rect 30716 43762 30772 44044
rect 30716 43710 30718 43762
rect 30770 43710 30772 43762
rect 30716 43698 30772 43710
rect 30268 43426 30324 43438
rect 30268 43374 30270 43426
rect 30322 43374 30324 43426
rect 30268 43204 30324 43374
rect 30268 43138 30324 43148
rect 30380 42868 30436 42878
rect 30156 42866 30436 42868
rect 30156 42814 30382 42866
rect 30434 42814 30436 42866
rect 30156 42812 30436 42814
rect 29932 42802 29988 42812
rect 30380 42802 30436 42812
rect 29596 42130 29652 42140
rect 29372 41918 29374 41970
rect 29426 41918 29428 41970
rect 28476 41858 28532 41870
rect 28476 41806 28478 41858
rect 28530 41806 28532 41858
rect 28476 41524 28532 41806
rect 28476 41458 28532 41468
rect 28028 41298 28196 41300
rect 28028 41246 28030 41298
rect 28082 41246 28196 41298
rect 28028 41244 28196 41246
rect 28028 41234 28084 41244
rect 29372 38948 29428 41918
rect 30940 41860 30996 45724
rect 31164 45714 31220 45724
rect 31052 45556 31108 45566
rect 31052 45332 31108 45500
rect 31164 45332 31220 45342
rect 31052 45330 31220 45332
rect 31052 45278 31166 45330
rect 31218 45278 31220 45330
rect 31052 45276 31220 45278
rect 31164 43762 31220 45276
rect 31164 43710 31166 43762
rect 31218 43710 31220 43762
rect 31164 43698 31220 43710
rect 31276 44098 31332 44110
rect 31276 44046 31278 44098
rect 31330 44046 31332 44098
rect 31276 43428 31332 44046
rect 31388 43652 31444 45838
rect 31948 45892 32004 45902
rect 31948 45798 32004 45836
rect 33180 45892 33236 47068
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 33852 46004 33908 46014
rect 35644 46004 35700 49200
rect 35756 46004 35812 46014
rect 35644 46002 35812 46004
rect 35644 45950 35758 46002
rect 35810 45950 35812 46002
rect 35644 45948 35812 45950
rect 33852 45910 33908 45948
rect 35756 45938 35812 45948
rect 33180 45890 33572 45892
rect 33180 45838 33182 45890
rect 33234 45838 33572 45890
rect 33180 45836 33572 45838
rect 33180 45826 33236 45836
rect 31724 45444 31780 45454
rect 31612 45220 31668 45230
rect 31612 45126 31668 45164
rect 31724 44434 31780 45388
rect 33516 45330 33572 45836
rect 35084 45890 35140 45902
rect 35084 45838 35086 45890
rect 35138 45838 35140 45890
rect 33516 45278 33518 45330
rect 33570 45278 33572 45330
rect 33516 45266 33572 45278
rect 34748 45332 34804 45342
rect 34748 45238 34804 45276
rect 35084 45332 35140 45838
rect 37660 45780 37716 49200
rect 37884 45780 37940 45790
rect 37660 45778 37940 45780
rect 37660 45726 37886 45778
rect 37938 45726 37940 45778
rect 37660 45724 37940 45726
rect 39676 45780 39732 49200
rect 42476 46452 42532 46462
rect 42476 46004 42532 46396
rect 43036 46004 43092 49200
rect 42476 46002 42980 46004
rect 42476 45950 42478 46002
rect 42530 45950 42980 46002
rect 42476 45948 42980 45950
rect 42476 45938 42532 45948
rect 42924 45890 42980 45948
rect 43036 45938 43092 45948
rect 43708 46004 43764 46014
rect 43708 45910 43764 45948
rect 42924 45838 42926 45890
rect 42978 45838 42980 45890
rect 42924 45826 42980 45838
rect 39900 45780 39956 45790
rect 39676 45778 39956 45780
rect 39676 45726 39902 45778
rect 39954 45726 39956 45778
rect 39676 45724 39956 45726
rect 37884 45714 37940 45724
rect 39900 45714 39956 45724
rect 48076 45780 48132 45790
rect 48412 45780 48468 49200
rect 48076 45778 48468 45780
rect 48076 45726 48078 45778
rect 48130 45726 48468 45778
rect 48076 45724 48468 45726
rect 48076 45714 48132 45724
rect 35084 45266 35140 45276
rect 32508 45108 32564 45118
rect 32508 45014 32564 45052
rect 31724 44382 31726 44434
rect 31778 44382 31780 44434
rect 31724 44370 31780 44382
rect 32060 44994 32116 45006
rect 32060 44942 32062 44994
rect 32114 44942 32116 44994
rect 31612 43652 31668 43662
rect 31388 43650 31668 43652
rect 31388 43598 31614 43650
rect 31666 43598 31668 43650
rect 31388 43596 31668 43598
rect 31612 43586 31668 43596
rect 32060 43652 32116 44942
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 32172 44436 32228 44446
rect 32172 44342 32228 44380
rect 32060 43586 32116 43596
rect 32620 44098 32676 44110
rect 32620 44046 32622 44098
rect 32674 44046 32676 44098
rect 31276 43362 31332 43372
rect 30940 41794 30996 41804
rect 32620 40628 32676 44046
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 32620 40562 32676 40572
rect 48076 40514 48132 40526
rect 48076 40462 48078 40514
rect 48130 40462 48132 40514
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 48076 39732 48132 40462
rect 48076 39666 48132 39676
rect 29372 38882 29428 38892
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 48076 37826 48132 37838
rect 48076 37774 48078 37826
rect 48130 37774 48132 37826
rect 48076 37716 48132 37774
rect 48076 37650 48132 37660
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 27916 36754 27972 36764
rect 27468 36530 27524 36540
rect 26796 35746 26852 35756
rect 48076 36258 48132 36270
rect 48076 36206 48078 36258
rect 48130 36206 48132 36258
rect 48076 35700 48132 36206
rect 48076 35634 48132 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 26236 35186 26292 35196
rect 21868 34962 21924 34972
rect 48076 34690 48132 34702
rect 48076 34638 48078 34690
rect 48130 34638 48132 34690
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 48076 34356 48132 34638
rect 48076 34290 48132 34300
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 19628 33506 19684 33516
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 48076 32674 48132 32686
rect 48076 32622 48078 32674
rect 48130 32622 48132 32674
rect 48076 32340 48132 32622
rect 48076 32274 48132 32284
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 48076 31554 48132 31566
rect 48076 31502 48078 31554
rect 48130 31502 48132 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 48076 30996 48132 31502
rect 48076 30930 48132 30940
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 48076 29538 48132 29550
rect 48076 29486 48078 29538
rect 48130 29486 48132 29538
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 48076 28980 48132 29486
rect 48076 28914 48132 28924
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 48076 26852 48132 26862
rect 48076 26758 48132 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 48076 23714 48132 23726
rect 48076 23662 48078 23714
rect 48130 23662 48132 23714
rect 48076 23604 48132 23662
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 48076 23538 48132 23548
rect 19836 23482 20100 23492
rect 11228 23314 11284 23324
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 48076 22146 48132 22158
rect 48076 22094 48078 22146
rect 48130 22094 48132 22146
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 48076 21588 48132 22094
rect 48076 21522 48132 21532
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 48076 18564 48132 18574
rect 48076 18470 48132 18508
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 48076 17442 48132 17454
rect 48076 17390 48078 17442
rect 48130 17390 48132 17442
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 48076 16884 48132 17390
rect 48076 16818 48132 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 48076 12852 48132 12862
rect 48076 12758 48132 12796
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 48076 12290 48132 12302
rect 48076 12238 48078 12290
rect 48130 12238 48132 12290
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 48076 11508 48132 12238
rect 48076 11442 48132 11452
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 48076 9602 48132 9614
rect 48076 9550 48078 9602
rect 48130 9550 48132 9602
rect 48076 9492 48132 9550
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 48076 9426 48132 9436
rect 19836 9370 20100 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 48076 8034 48132 8046
rect 48076 7982 48078 8034
rect 48130 7982 48132 8034
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 48076 7476 48132 7982
rect 48076 7410 48132 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 48076 6466 48132 6478
rect 48076 6414 48078 6466
rect 48130 6414 48132 6466
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 48076 6132 48132 6414
rect 48076 6066 48132 6076
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 5852 3602 5908 3612
rect 3052 3502 3054 3554
rect 3106 3502 3108 3554
rect 3052 3490 3108 3502
rect 3612 3332 3668 3342
rect 2492 2258 2548 2268
rect 3388 3330 3668 3332
rect 3388 3278 3614 3330
rect 3666 3278 3668 3330
rect 3388 3276 3668 3278
rect 3388 800 3444 3276
rect 3612 3266 3668 3276
rect 4732 3332 4788 3342
rect 4732 800 4788 3276
rect 5740 3332 5796 3342
rect 5740 3238 5796 3276
rect 9660 3330 9716 3342
rect 14364 3332 14420 3342
rect 15708 3332 15764 3342
rect 17724 3332 17780 3342
rect 9660 3278 9662 3330
rect 9714 3278 9716 3330
rect 8764 1762 8820 1774
rect 8764 1710 8766 1762
rect 8818 1710 8820 1762
rect 8764 800 8820 1710
rect 9660 1762 9716 3278
rect 9660 1710 9662 1762
rect 9714 1710 9716 1762
rect 9660 1698 9716 1710
rect 14140 3330 14420 3332
rect 14140 3278 14366 3330
rect 14418 3278 14420 3330
rect 14140 3276 14420 3278
rect 14140 800 14196 3276
rect 14364 3266 14420 3276
rect 15484 3330 15764 3332
rect 15484 3278 15710 3330
rect 15762 3278 15764 3330
rect 15484 3276 15764 3278
rect 15484 800 15540 3276
rect 15708 3266 15764 3276
rect 17500 3330 17780 3332
rect 17500 3278 17726 3330
rect 17778 3278 17780 3330
rect 17500 3276 17780 3278
rect 17500 800 17556 3276
rect 17724 3266 17780 3276
rect 21420 3330 21476 3342
rect 23100 3332 23156 3342
rect 26460 3332 26516 3342
rect 21420 3278 21422 3330
rect 21474 3278 21476 3330
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 1762 20916 1774
rect 20860 1710 20862 1762
rect 20914 1710 20916 1762
rect 20860 800 20916 1710
rect 21420 1762 21476 3278
rect 21420 1710 21422 1762
rect 21474 1710 21476 1762
rect 21420 1698 21476 1710
rect 22876 3330 23156 3332
rect 22876 3278 23102 3330
rect 23154 3278 23156 3330
rect 22876 3276 23156 3278
rect 22876 800 22932 3276
rect 23100 3266 23156 3276
rect 26236 3330 26516 3332
rect 26236 3278 26462 3330
rect 26514 3278 26516 3330
rect 26236 3276 26516 3278
rect 26236 800 26292 3276
rect 26460 3266 26516 3276
rect 28252 3332 28308 3342
rect 28252 800 28308 3276
rect 29260 3332 29316 3342
rect 31836 3332 31892 3342
rect 35196 3332 35252 3342
rect 38556 3332 38612 3342
rect 29260 3238 29316 3276
rect 31612 3330 31892 3332
rect 31612 3278 31838 3330
rect 31890 3278 31892 3330
rect 31612 3276 31892 3278
rect 31612 800 31668 3276
rect 31836 3266 31892 3276
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 38332 3330 38612 3332
rect 38332 3278 38558 3330
rect 38610 3278 38612 3330
rect 38332 3276 38612 3278
rect 38332 800 38388 3276
rect 38556 3266 38612 3276
rect 41020 3330 41076 3342
rect 42588 3332 42644 3342
rect 43932 3332 43988 3342
rect 45948 3332 46004 3342
rect 41020 3278 41022 3330
rect 41074 3278 41076 3330
rect 40348 1874 40404 1886
rect 40348 1822 40350 1874
rect 40402 1822 40404 1874
rect 40348 800 40404 1822
rect 41020 1874 41076 3278
rect 41020 1822 41022 1874
rect 41074 1822 41076 1874
rect 41020 1810 41076 1822
rect 42364 3330 42644 3332
rect 42364 3278 42590 3330
rect 42642 3278 42644 3330
rect 42364 3276 42644 3278
rect 42364 800 42420 3276
rect 42588 3266 42644 3276
rect 43708 3330 43988 3332
rect 43708 3278 43934 3330
rect 43986 3278 43988 3330
rect 43708 3276 43988 3278
rect 43708 800 43764 3276
rect 43932 3266 43988 3276
rect 45724 3330 46004 3332
rect 45724 3278 45950 3330
rect 46002 3278 46004 3330
rect 45724 3276 46004 3278
rect 45724 800 45780 3276
rect 45948 3266 46004 3276
rect 47404 3330 47460 3342
rect 47404 3278 47406 3330
rect 47458 3278 47460 3330
rect 47404 2100 47460 3278
rect 47404 2034 47460 2044
rect 48076 3330 48132 3342
rect 48076 3278 48078 3330
rect 48130 3278 48132 3330
rect 0 200 112 800
rect 1344 200 1456 800
rect 3360 200 3472 800
rect 4704 200 4816 800
rect 6720 200 6832 800
rect 8736 200 8848 800
rect 10080 200 10192 800
rect 12096 200 12208 800
rect 14112 200 14224 800
rect 15456 200 15568 800
rect 17472 200 17584 800
rect 18816 200 18928 800
rect 20832 200 20944 800
rect 22848 200 22960 800
rect 24192 200 24304 800
rect 26208 200 26320 800
rect 28224 200 28336 800
rect 29568 200 29680 800
rect 31584 200 31696 800
rect 33600 200 33712 800
rect 34944 200 35056 800
rect 36960 200 37072 800
rect 38304 200 38416 800
rect 40320 200 40432 800
rect 42336 200 42448 800
rect 43680 200 43792 800
rect 45696 200 45808 800
rect 47712 200 47824 800
rect 48076 756 48132 3278
rect 48076 690 48132 700
rect 49056 200 49168 800
<< via2 >>
rect 3388 49084 3444 49140
rect 2492 45724 2548 45780
rect 1820 45666 1876 45668
rect 1820 45614 1822 45666
rect 1822 45614 1874 45666
rect 1874 45614 1876 45666
rect 1820 45612 1876 45614
rect 3052 46396 3108 46452
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 6860 46060 6916 46116
rect 4956 45890 5012 45892
rect 4956 45838 4958 45890
rect 4958 45838 5010 45890
rect 5010 45838 5012 45890
rect 4956 45836 5012 45838
rect 3500 45612 3556 45668
rect 3164 45330 3220 45332
rect 3164 45278 3166 45330
rect 3166 45278 3218 45330
rect 3218 45278 3220 45330
rect 3164 45276 3220 45278
rect 4284 45612 4340 45668
rect 4172 45500 4228 45556
rect 3724 44434 3780 44436
rect 3724 44382 3726 44434
rect 3726 44382 3778 44434
rect 3778 44382 3780 44434
rect 3724 44380 3780 44382
rect 2156 43708 2212 43764
rect 4284 45052 4340 45108
rect 4060 43820 4116 43876
rect 5516 45612 5572 45668
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4620 44098 4676 44100
rect 4620 44046 4622 44098
rect 4622 44046 4674 44098
rect 4674 44046 4676 44098
rect 4620 44044 4676 44046
rect 4956 44994 5012 44996
rect 4956 44942 4958 44994
rect 4958 44942 5010 44994
rect 5010 44942 5012 44994
rect 4956 44940 5012 44942
rect 3500 43426 3556 43428
rect 3500 43374 3502 43426
rect 3502 43374 3554 43426
rect 3554 43374 3556 43426
rect 3500 43372 3556 43374
rect 3948 42812 4004 42868
rect 1820 42364 1876 42420
rect 4844 43762 4900 43764
rect 4844 43710 4846 43762
rect 4846 43710 4898 43762
rect 4898 43710 4900 43762
rect 4844 43708 4900 43710
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4508 42866 4564 42868
rect 4508 42814 4510 42866
rect 4510 42814 4562 42866
rect 4562 42814 4564 42866
rect 4508 42812 4564 42814
rect 4284 42140 4340 42196
rect 5068 43932 5124 43988
rect 5180 43820 5236 43876
rect 5068 43596 5124 43652
rect 5180 43484 5236 43540
rect 5740 45388 5796 45444
rect 5404 43372 5460 43428
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4956 41580 5012 41636
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5852 44268 5908 44324
rect 5628 42194 5684 42196
rect 5628 42142 5630 42194
rect 5630 42142 5682 42194
rect 5682 42142 5684 42194
rect 5628 42140 5684 42142
rect 5628 41020 5684 41076
rect 5404 39788 5460 39844
rect 6188 45106 6244 45108
rect 6188 45054 6190 45106
rect 6190 45054 6242 45106
rect 6242 45054 6244 45106
rect 6188 45052 6244 45054
rect 6524 44322 6580 44324
rect 6524 44270 6526 44322
rect 6526 44270 6578 44322
rect 6578 44270 6580 44322
rect 6524 44268 6580 44270
rect 6748 43820 6804 43876
rect 6076 43596 6132 43652
rect 6188 42140 6244 42196
rect 6636 42924 6692 42980
rect 6300 41916 6356 41972
rect 6076 41692 6132 41748
rect 5964 39004 6020 39060
rect 6412 41298 6468 41300
rect 6412 41246 6414 41298
rect 6414 41246 6466 41298
rect 6466 41246 6468 41298
rect 6412 41244 6468 41246
rect 1820 38332 1876 38388
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 6636 40124 6692 40180
rect 7308 44210 7364 44212
rect 7308 44158 7310 44210
rect 7310 44158 7362 44210
rect 7362 44158 7364 44210
rect 7308 44156 7364 44158
rect 7980 45948 8036 46004
rect 7420 43820 7476 43876
rect 7756 45164 7812 45220
rect 7308 43426 7364 43428
rect 7308 43374 7310 43426
rect 7310 43374 7362 43426
rect 7362 43374 7364 43426
rect 7308 43372 7364 43374
rect 7308 42812 7364 42868
rect 7084 42754 7140 42756
rect 7084 42702 7086 42754
rect 7086 42702 7138 42754
rect 7138 42702 7140 42754
rect 7084 42700 7140 42702
rect 7644 42812 7700 42868
rect 7084 41858 7140 41860
rect 7084 41806 7086 41858
rect 7086 41806 7138 41858
rect 7138 41806 7140 41858
rect 7084 41804 7140 41806
rect 7532 42028 7588 42084
rect 7420 41692 7476 41748
rect 7308 41468 7364 41524
rect 7868 44492 7924 44548
rect 7868 43708 7924 43764
rect 8092 45778 8148 45780
rect 8092 45726 8094 45778
rect 8094 45726 8146 45778
rect 8146 45726 8148 45778
rect 8092 45724 8148 45726
rect 11340 48188 11396 48244
rect 10668 48076 10724 48132
rect 9996 47740 10052 47796
rect 9548 45724 9604 45780
rect 8764 45052 8820 45108
rect 8988 45164 9044 45220
rect 8988 43708 9044 43764
rect 8876 43650 8932 43652
rect 8876 43598 8878 43650
rect 8878 43598 8930 43650
rect 8930 43598 8932 43650
rect 8876 43596 8932 43598
rect 8764 43484 8820 43540
rect 8540 43372 8596 43428
rect 7980 42812 8036 42868
rect 8204 42700 8260 42756
rect 8092 42530 8148 42532
rect 8092 42478 8094 42530
rect 8094 42478 8146 42530
rect 8146 42478 8148 42530
rect 8092 42476 8148 42478
rect 7980 41356 8036 41412
rect 8092 41580 8148 41636
rect 8428 43036 8484 43092
rect 8204 40402 8260 40404
rect 8204 40350 8206 40402
rect 8206 40350 8258 40402
rect 8258 40350 8260 40402
rect 8204 40348 8260 40350
rect 8316 40012 8372 40068
rect 7196 39340 7252 39396
rect 6748 38892 6804 38948
rect 6412 37884 6468 37940
rect 8876 43426 8932 43428
rect 8876 43374 8878 43426
rect 8878 43374 8930 43426
rect 8930 43374 8932 43426
rect 8876 43372 8932 43374
rect 8652 42642 8708 42644
rect 8652 42590 8654 42642
rect 8654 42590 8706 42642
rect 8706 42590 8708 42642
rect 8652 42588 8708 42590
rect 8764 42140 8820 42196
rect 8652 41580 8708 41636
rect 10668 45500 10724 45556
rect 10892 47628 10948 47684
rect 9996 45276 10052 45332
rect 9548 44940 9604 44996
rect 9100 41186 9156 41188
rect 9100 41134 9102 41186
rect 9102 41134 9154 41186
rect 9154 41134 9156 41186
rect 9100 41132 9156 41134
rect 9324 43036 9380 43092
rect 9660 44828 9716 44884
rect 9660 43762 9716 43764
rect 9660 43710 9662 43762
rect 9662 43710 9714 43762
rect 9714 43710 9716 43762
rect 9660 43708 9716 43710
rect 10108 45106 10164 45108
rect 10108 45054 10110 45106
rect 10110 45054 10162 45106
rect 10162 45054 10164 45106
rect 10108 45052 10164 45054
rect 10108 43708 10164 43764
rect 9212 40460 9268 40516
rect 9436 42700 9492 42756
rect 9884 42700 9940 42756
rect 9996 42588 10052 42644
rect 9996 42364 10052 42420
rect 9996 41804 10052 41860
rect 9660 41692 9716 41748
rect 9548 41298 9604 41300
rect 9548 41246 9550 41298
rect 9550 41246 9602 41298
rect 9602 41246 9604 41298
rect 9548 41244 9604 41246
rect 9996 41020 10052 41076
rect 9660 40572 9716 40628
rect 10332 43708 10388 43764
rect 10444 44268 10500 44324
rect 10220 42812 10276 42868
rect 10220 41970 10276 41972
rect 10220 41918 10222 41970
rect 10222 41918 10274 41970
rect 10274 41918 10276 41970
rect 10220 41916 10276 41918
rect 10668 43932 10724 43988
rect 10556 43036 10612 43092
rect 10332 41468 10388 41524
rect 10220 40626 10276 40628
rect 10220 40574 10222 40626
rect 10222 40574 10274 40626
rect 10274 40574 10276 40626
rect 10220 40572 10276 40574
rect 10780 42476 10836 42532
rect 11116 45106 11172 45108
rect 11116 45054 11118 45106
rect 11118 45054 11170 45106
rect 11170 45054 11172 45106
rect 11116 45052 11172 45054
rect 11004 44716 11060 44772
rect 11228 44492 11284 44548
rect 11004 44380 11060 44436
rect 10892 42194 10948 42196
rect 10892 42142 10894 42194
rect 10894 42142 10946 42194
rect 10946 42142 10948 42194
rect 10892 42140 10948 42142
rect 11228 44156 11284 44212
rect 11452 47628 11508 47684
rect 11452 44994 11508 44996
rect 11452 44942 11454 44994
rect 11454 44942 11506 44994
rect 11506 44942 11508 44994
rect 11452 44940 11508 44942
rect 11676 44882 11732 44884
rect 11676 44830 11678 44882
rect 11678 44830 11730 44882
rect 11730 44830 11732 44882
rect 11676 44828 11732 44830
rect 11564 44492 11620 44548
rect 11452 44156 11508 44212
rect 11452 43932 11508 43988
rect 11340 42924 11396 42980
rect 11564 42924 11620 42980
rect 11452 42476 11508 42532
rect 11340 42028 11396 42084
rect 11340 41468 11396 41524
rect 11564 42364 11620 42420
rect 11340 40908 11396 40964
rect 11452 41020 11508 41076
rect 11340 40514 11396 40516
rect 11340 40462 11342 40514
rect 11342 40462 11394 40514
rect 11394 40462 11396 40514
rect 11340 40460 11396 40462
rect 10108 40348 10164 40404
rect 10556 40348 10612 40404
rect 9548 39730 9604 39732
rect 9548 39678 9550 39730
rect 9550 39678 9602 39730
rect 9602 39678 9604 39730
rect 9548 39676 9604 39678
rect 9996 39730 10052 39732
rect 9996 39678 9998 39730
rect 9998 39678 10050 39730
rect 10050 39678 10052 39730
rect 9996 39676 10052 39678
rect 9436 39116 9492 39172
rect 10556 39730 10612 39732
rect 10556 39678 10558 39730
rect 10558 39678 10610 39730
rect 10610 39678 10612 39730
rect 10556 39676 10612 39678
rect 10108 38556 10164 38612
rect 10444 39116 10500 39172
rect 10892 38556 10948 38612
rect 10556 38162 10612 38164
rect 10556 38110 10558 38162
rect 10558 38110 10610 38162
rect 10610 38110 10612 38162
rect 10556 38108 10612 38110
rect 10444 37324 10500 37380
rect 8540 37212 8596 37268
rect 1820 36988 1876 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 11340 39058 11396 39060
rect 11340 39006 11342 39058
rect 11342 39006 11394 39058
rect 11394 39006 11396 39058
rect 11340 39004 11396 39006
rect 16716 47964 16772 48020
rect 14028 47852 14084 47908
rect 12796 46508 12852 46564
rect 12236 46396 12292 46452
rect 12124 45724 12180 45780
rect 12124 45388 12180 45444
rect 13580 45890 13636 45892
rect 13580 45838 13582 45890
rect 13582 45838 13634 45890
rect 13634 45838 13636 45890
rect 13580 45836 13636 45838
rect 12572 43372 12628 43428
rect 12124 42364 12180 42420
rect 12908 42476 12964 42532
rect 12572 42028 12628 42084
rect 11676 41132 11732 41188
rect 11564 37660 11620 37716
rect 11452 37436 11508 37492
rect 11116 36764 11172 36820
rect 5852 36092 5908 36148
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1820 34972 1876 35028
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 1820 32956 1876 33012
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1820 29596 1876 29652
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 1820 28252 1876 28308
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 1820 26236 1876 26292
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1820 24220 1876 24276
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 3052 23324 3108 23380
rect 3500 23378 3556 23380
rect 3500 23326 3502 23378
rect 3502 23326 3554 23378
rect 3554 23326 3556 23378
rect 3500 23324 3556 23326
rect 2044 22876 2100 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1820 20860 1876 20916
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 1820 18844 1876 18900
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1820 17554 1876 17556
rect 1820 17502 1822 17554
rect 1822 17502 1874 17554
rect 1874 17502 1876 17554
rect 1820 17500 1876 17502
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1820 15484 1876 15540
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 1820 14140 1876 14196
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 1820 10108 1876 10164
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 1820 8764 1876 8820
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 1820 6748 1876 6804
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 1372 3500 1428 3556
rect 28 2268 84 2324
rect 2156 3554 2212 3556
rect 2156 3502 2158 3554
rect 2158 3502 2210 3554
rect 2210 3502 2212 3554
rect 2156 3500 2212 3502
rect 1820 3388 1876 3444
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 3052 3612 3108 3668
rect 4284 3666 4340 3668
rect 4284 3614 4286 3666
rect 4286 3614 4338 3666
rect 4338 3614 4340 3666
rect 4284 3612 4340 3614
rect 11228 35532 11284 35588
rect 11900 39900 11956 39956
rect 12124 40348 12180 40404
rect 12348 40012 12404 40068
rect 12908 41356 12964 41412
rect 13692 43484 13748 43540
rect 13468 43426 13524 43428
rect 13468 43374 13470 43426
rect 13470 43374 13522 43426
rect 13522 43374 13524 43426
rect 13468 43372 13524 43374
rect 13692 43148 13748 43204
rect 15708 47516 15764 47572
rect 14476 45836 14532 45892
rect 14140 44098 14196 44100
rect 14140 44046 14142 44098
rect 14142 44046 14194 44098
rect 14194 44046 14196 44098
rect 14140 44044 14196 44046
rect 14028 43484 14084 43540
rect 13916 42978 13972 42980
rect 13916 42926 13918 42978
rect 13918 42926 13970 42978
rect 13970 42926 13972 42978
rect 13916 42924 13972 42926
rect 13916 42364 13972 42420
rect 13692 41692 13748 41748
rect 13020 40124 13076 40180
rect 13244 41356 13300 41412
rect 12572 39900 12628 39956
rect 12796 39564 12852 39620
rect 12012 38556 12068 38612
rect 12908 39506 12964 39508
rect 12908 39454 12910 39506
rect 12910 39454 12962 39506
rect 12962 39454 12964 39506
rect 12908 39452 12964 39454
rect 12684 38108 12740 38164
rect 13692 41132 13748 41188
rect 13804 42252 13860 42308
rect 13692 40460 13748 40516
rect 14364 43036 14420 43092
rect 14924 45276 14980 45332
rect 14588 45106 14644 45108
rect 14588 45054 14590 45106
rect 14590 45054 14642 45106
rect 14642 45054 14644 45106
rect 14588 45052 14644 45054
rect 14588 44828 14644 44884
rect 14364 42754 14420 42756
rect 14364 42702 14366 42754
rect 14366 42702 14418 42754
rect 14418 42702 14420 42754
rect 14364 42700 14420 42702
rect 14364 42140 14420 42196
rect 14588 41804 14644 41860
rect 15372 45276 15428 45332
rect 15148 44380 15204 44436
rect 14924 42476 14980 42532
rect 14476 41692 14532 41748
rect 14924 41356 14980 41412
rect 15036 42588 15092 42644
rect 14028 39676 14084 39732
rect 14140 40908 14196 40964
rect 14924 40962 14980 40964
rect 14924 40910 14926 40962
rect 14926 40910 14978 40962
rect 14978 40910 14980 40962
rect 14924 40908 14980 40910
rect 14812 40796 14868 40852
rect 14364 40572 14420 40628
rect 14924 40402 14980 40404
rect 14924 40350 14926 40402
rect 14926 40350 14978 40402
rect 14978 40350 14980 40402
rect 14924 40348 14980 40350
rect 14364 40236 14420 40292
rect 15596 44380 15652 44436
rect 16604 47404 16660 47460
rect 16044 47292 16100 47348
rect 15932 45890 15988 45892
rect 15932 45838 15934 45890
rect 15934 45838 15986 45890
rect 15986 45838 15988 45890
rect 15932 45836 15988 45838
rect 15820 45164 15876 45220
rect 15932 44994 15988 44996
rect 15932 44942 15934 44994
rect 15934 44942 15986 44994
rect 15986 44942 15988 44994
rect 15932 44940 15988 44942
rect 15820 44156 15876 44212
rect 15260 42924 15316 42980
rect 15148 41580 15204 41636
rect 15036 39676 15092 39732
rect 15148 41356 15204 41412
rect 14028 39004 14084 39060
rect 13020 38162 13076 38164
rect 13020 38110 13022 38162
rect 13022 38110 13074 38162
rect 13074 38110 13076 38162
rect 13020 38108 13076 38110
rect 12684 37100 12740 37156
rect 14252 39340 14308 39396
rect 14252 38780 14308 38836
rect 15484 42140 15540 42196
rect 15708 43260 15764 43316
rect 15708 43036 15764 43092
rect 15708 42812 15764 42868
rect 15596 41580 15652 41636
rect 15484 41020 15540 41076
rect 15820 41804 15876 41860
rect 16268 46172 16324 46228
rect 16380 45612 16436 45668
rect 16492 45276 16548 45332
rect 16380 45106 16436 45108
rect 16380 45054 16382 45106
rect 16382 45054 16434 45106
rect 16434 45054 16436 45106
rect 16380 45052 16436 45054
rect 16156 44156 16212 44212
rect 16492 44716 16548 44772
rect 16268 44098 16324 44100
rect 16268 44046 16270 44098
rect 16270 44046 16322 44098
rect 16322 44046 16324 44098
rect 16268 44044 16324 44046
rect 16156 43036 16212 43092
rect 16044 42812 16100 42868
rect 16044 42364 16100 42420
rect 16268 42028 16324 42084
rect 16156 41580 16212 41636
rect 15820 41132 15876 41188
rect 15708 40572 15764 40628
rect 15820 40684 15876 40740
rect 15148 39564 15204 39620
rect 15372 40124 15428 40180
rect 14812 39116 14868 39172
rect 14812 37938 14868 37940
rect 14812 37886 14814 37938
rect 14814 37886 14866 37938
rect 14866 37886 14868 37938
rect 14812 37884 14868 37886
rect 14588 37490 14644 37492
rect 14588 37438 14590 37490
rect 14590 37438 14642 37490
rect 14642 37438 14644 37490
rect 14588 37436 14644 37438
rect 14924 37154 14980 37156
rect 14924 37102 14926 37154
rect 14926 37102 14978 37154
rect 14978 37102 14980 37154
rect 14924 37100 14980 37102
rect 14364 36652 14420 36708
rect 13916 36540 13972 36596
rect 13692 36204 13748 36260
rect 12124 36092 12180 36148
rect 15260 36876 15316 36932
rect 15260 36652 15316 36708
rect 15036 36540 15092 36596
rect 15820 40124 15876 40180
rect 15596 40012 15652 40068
rect 15596 39676 15652 39732
rect 15708 39900 15764 39956
rect 15484 39116 15540 39172
rect 15596 39228 15652 39284
rect 15596 38108 15652 38164
rect 15484 37436 15540 37492
rect 15484 37266 15540 37268
rect 15484 37214 15486 37266
rect 15486 37214 15538 37266
rect 15538 37214 15540 37266
rect 15484 37212 15540 37214
rect 15148 36428 15204 36484
rect 15596 36428 15652 36484
rect 14700 35980 14756 36036
rect 15260 35980 15316 36036
rect 11788 35532 11844 35588
rect 15820 39340 15876 39396
rect 16156 41132 16212 41188
rect 16380 41804 16436 41860
rect 16380 41580 16436 41636
rect 16380 41356 16436 41412
rect 16268 40684 16324 40740
rect 16380 41020 16436 41076
rect 17836 45724 17892 45780
rect 17500 45666 17556 45668
rect 17500 45614 17502 45666
rect 17502 45614 17554 45666
rect 17554 45614 17556 45666
rect 17500 45612 17556 45614
rect 16716 45164 16772 45220
rect 16828 44322 16884 44324
rect 16828 44270 16830 44322
rect 16830 44270 16882 44322
rect 16882 44270 16884 44322
rect 16828 44268 16884 44270
rect 16828 43708 16884 43764
rect 17388 44156 17444 44212
rect 16604 43260 16660 43316
rect 16604 42476 16660 42532
rect 16604 41468 16660 41524
rect 16716 41244 16772 41300
rect 16828 43260 16884 43316
rect 16828 42028 16884 42084
rect 16604 40572 16660 40628
rect 16380 39452 16436 39508
rect 16940 40684 16996 40740
rect 17052 41804 17108 41860
rect 16940 40514 16996 40516
rect 16940 40462 16942 40514
rect 16942 40462 16994 40514
rect 16994 40462 16996 40514
rect 16940 40460 16996 40462
rect 16828 39340 16884 39396
rect 16156 39228 16212 39284
rect 16044 39004 16100 39060
rect 16716 39004 16772 39060
rect 16044 38780 16100 38836
rect 16156 38892 16212 38948
rect 16716 37996 16772 38052
rect 15932 37154 15988 37156
rect 15932 37102 15934 37154
rect 15934 37102 15986 37154
rect 15986 37102 15988 37154
rect 15932 37100 15988 37102
rect 16044 37042 16100 37044
rect 16044 36990 16046 37042
rect 16046 36990 16098 37042
rect 16098 36990 16100 37042
rect 16044 36988 16100 36990
rect 15932 36876 15988 36932
rect 16156 36652 16212 36708
rect 16604 37266 16660 37268
rect 16604 37214 16606 37266
rect 16606 37214 16658 37266
rect 16658 37214 16660 37266
rect 16604 37212 16660 37214
rect 16716 36988 16772 37044
rect 16828 36652 16884 36708
rect 17388 39900 17444 39956
rect 17276 39788 17332 39844
rect 17164 39618 17220 39620
rect 17164 39566 17166 39618
rect 17166 39566 17218 39618
rect 17218 39566 17220 39618
rect 17164 39564 17220 39566
rect 17052 38834 17108 38836
rect 17052 38782 17054 38834
rect 17054 38782 17106 38834
rect 17106 38782 17108 38834
rect 17052 38780 17108 38782
rect 16716 36482 16772 36484
rect 16716 36430 16718 36482
rect 16718 36430 16770 36482
rect 16770 36430 16772 36482
rect 16716 36428 16772 36430
rect 17724 43148 17780 43204
rect 19404 46732 19460 46788
rect 18956 45612 19012 45668
rect 18396 45388 18452 45444
rect 17724 42028 17780 42084
rect 18396 45218 18452 45220
rect 18396 45166 18398 45218
rect 18398 45166 18450 45218
rect 18450 45166 18452 45218
rect 18396 45164 18452 45166
rect 18172 43932 18228 43988
rect 18060 42252 18116 42308
rect 18172 43148 18228 43204
rect 17948 41804 18004 41860
rect 17836 41468 17892 41524
rect 18060 41692 18116 41748
rect 17724 41356 17780 41412
rect 17948 40236 18004 40292
rect 17388 39676 17444 39732
rect 17276 38108 17332 38164
rect 17500 39452 17556 39508
rect 17948 39452 18004 39508
rect 17612 39116 17668 39172
rect 17836 38946 17892 38948
rect 17836 38894 17838 38946
rect 17838 38894 17890 38946
rect 17890 38894 17892 38946
rect 17836 38892 17892 38894
rect 17724 38834 17780 38836
rect 17724 38782 17726 38834
rect 17726 38782 17778 38834
rect 17778 38782 17780 38834
rect 17724 38780 17780 38782
rect 17948 37772 18004 37828
rect 19180 43932 19236 43988
rect 18284 42028 18340 42084
rect 18508 41916 18564 41972
rect 18620 42812 18676 42868
rect 18172 40348 18228 40404
rect 18508 39900 18564 39956
rect 18396 39340 18452 39396
rect 18508 38668 18564 38724
rect 19068 41804 19124 41860
rect 18732 41298 18788 41300
rect 18732 41246 18734 41298
rect 18734 41246 18786 41298
rect 18786 41246 18788 41298
rect 18732 41244 18788 41246
rect 18956 40124 19012 40180
rect 18844 38834 18900 38836
rect 18844 38782 18846 38834
rect 18846 38782 18898 38834
rect 18898 38782 18900 38834
rect 18844 38780 18900 38782
rect 19292 39788 19348 39844
rect 19292 39058 19348 39060
rect 19292 39006 19294 39058
rect 19294 39006 19346 39058
rect 19346 39006 19348 39058
rect 19292 39004 19348 39006
rect 19180 38780 19236 38836
rect 19068 38668 19124 38724
rect 19964 45890 20020 45892
rect 19964 45838 19966 45890
rect 19966 45838 20018 45890
rect 20018 45838 20020 45890
rect 19964 45836 20020 45838
rect 19628 45500 19684 45556
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20300 47180 20356 47236
rect 20300 45948 20356 46004
rect 19628 44492 19684 44548
rect 20524 47068 20580 47124
rect 21084 45948 21140 46004
rect 20636 45276 20692 45332
rect 20972 45164 21028 45220
rect 20860 44716 20916 44772
rect 20860 44210 20916 44212
rect 20860 44158 20862 44210
rect 20862 44158 20914 44210
rect 20914 44158 20916 44210
rect 20860 44156 20916 44158
rect 20188 44044 20244 44100
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19628 43372 19684 43428
rect 20076 42812 20132 42868
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19964 42028 20020 42084
rect 19852 40908 19908 40964
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19852 40572 19908 40628
rect 20636 44098 20692 44100
rect 20636 44046 20638 44098
rect 20638 44046 20690 44098
rect 20690 44046 20692 44098
rect 20636 44044 20692 44046
rect 20636 43820 20692 43876
rect 20860 42924 20916 42980
rect 20748 42866 20804 42868
rect 20748 42814 20750 42866
rect 20750 42814 20802 42866
rect 20802 42814 20804 42866
rect 20748 42812 20804 42814
rect 20524 42140 20580 42196
rect 20636 42028 20692 42084
rect 20300 41580 20356 41636
rect 20412 41468 20468 41524
rect 20300 41132 20356 41188
rect 20300 40684 20356 40740
rect 20524 41356 20580 41412
rect 20860 42476 20916 42532
rect 20748 41804 20804 41860
rect 21420 45106 21476 45108
rect 21420 45054 21422 45106
rect 21422 45054 21474 45106
rect 21474 45054 21476 45106
rect 21420 45052 21476 45054
rect 21308 44716 21364 44772
rect 21196 43426 21252 43428
rect 21196 43374 21198 43426
rect 21198 43374 21250 43426
rect 21250 43374 21252 43426
rect 21196 43372 21252 43374
rect 24220 48188 24276 48244
rect 22092 45500 22148 45556
rect 25452 48076 25508 48132
rect 24892 46508 24948 46564
rect 24444 46396 24500 46452
rect 24668 46060 24724 46116
rect 24220 45388 24276 45444
rect 23772 45330 23828 45332
rect 23772 45278 23774 45330
rect 23774 45278 23826 45330
rect 23826 45278 23828 45330
rect 23772 45276 23828 45278
rect 24444 45500 24500 45556
rect 22316 44604 22372 44660
rect 21644 43484 21700 43540
rect 21980 43484 22036 43540
rect 21532 43372 21588 43428
rect 21196 42924 21252 42980
rect 20860 41468 20916 41524
rect 20636 41132 20692 41188
rect 20748 41020 20804 41076
rect 20412 40348 20468 40404
rect 20748 40348 20804 40404
rect 20300 39730 20356 39732
rect 20300 39678 20302 39730
rect 20302 39678 20354 39730
rect 20354 39678 20356 39730
rect 20300 39676 20356 39678
rect 20636 39564 20692 39620
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19964 38780 20020 38836
rect 19852 38722 19908 38724
rect 19852 38670 19854 38722
rect 19854 38670 19906 38722
rect 19906 38670 19908 38722
rect 19852 38668 19908 38670
rect 18284 37378 18340 37380
rect 18284 37326 18286 37378
rect 18286 37326 18338 37378
rect 18338 37326 18340 37378
rect 18284 37324 18340 37326
rect 17500 36764 17556 36820
rect 17612 36370 17668 36372
rect 17612 36318 17614 36370
rect 17614 36318 17666 36370
rect 17666 36318 17668 36370
rect 17612 36316 17668 36318
rect 18732 37772 18788 37828
rect 18396 36428 18452 36484
rect 18508 37436 18564 37492
rect 18508 37100 18564 37156
rect 18620 36316 18676 36372
rect 17276 36092 17332 36148
rect 18060 36092 18116 36148
rect 18284 36092 18340 36148
rect 18620 35922 18676 35924
rect 18620 35870 18622 35922
rect 18622 35870 18674 35922
rect 18674 35870 18676 35922
rect 18620 35868 18676 35870
rect 16604 35644 16660 35700
rect 15708 35196 15764 35252
rect 17948 35532 18004 35588
rect 17500 35026 17556 35028
rect 17500 34974 17502 35026
rect 17502 34974 17554 35026
rect 17554 34974 17556 35026
rect 17500 34972 17556 34974
rect 19180 38444 19236 38500
rect 18956 38220 19012 38276
rect 19180 37826 19236 37828
rect 19180 37774 19182 37826
rect 19182 37774 19234 37826
rect 19234 37774 19236 37826
rect 19180 37772 19236 37774
rect 19068 37660 19124 37716
rect 19292 37660 19348 37716
rect 19180 37548 19236 37604
rect 18956 36988 19012 37044
rect 19068 37100 19124 37156
rect 19180 36428 19236 36484
rect 19180 36092 19236 36148
rect 19404 37548 19460 37604
rect 19964 38556 20020 38612
rect 19628 38444 19684 38500
rect 19964 38332 20020 38388
rect 20412 38444 20468 38500
rect 20188 38332 20244 38388
rect 20076 38220 20132 38276
rect 20412 37938 20468 37940
rect 20412 37886 20414 37938
rect 20414 37886 20466 37938
rect 20466 37886 20468 37938
rect 20412 37884 20468 37886
rect 19628 37660 19684 37716
rect 20300 37772 20356 37828
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37436 20132 37492
rect 19740 37154 19796 37156
rect 19740 37102 19742 37154
rect 19742 37102 19794 37154
rect 19794 37102 19796 37154
rect 19740 37100 19796 37102
rect 19516 36988 19572 37044
rect 19964 36258 20020 36260
rect 19964 36206 19966 36258
rect 19966 36206 20018 36258
rect 20018 36206 20020 36258
rect 19964 36204 20020 36206
rect 20300 37154 20356 37156
rect 20300 37102 20302 37154
rect 20302 37102 20354 37154
rect 20354 37102 20356 37154
rect 20300 37100 20356 37102
rect 20524 37324 20580 37380
rect 20524 36988 20580 37044
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20972 40348 21028 40404
rect 20860 40012 20916 40068
rect 20860 38668 20916 38724
rect 20860 38332 20916 38388
rect 21196 41132 21252 41188
rect 21756 42140 21812 42196
rect 21084 38444 21140 38500
rect 20972 37436 21028 37492
rect 21308 39788 21364 39844
rect 21644 40796 21700 40852
rect 21756 40124 21812 40180
rect 21868 39788 21924 39844
rect 22092 41804 22148 41860
rect 22092 41074 22148 41076
rect 22092 41022 22094 41074
rect 22094 41022 22146 41074
rect 22146 41022 22148 41074
rect 22092 41020 22148 41022
rect 22428 44380 22484 44436
rect 22428 43932 22484 43988
rect 24444 44492 24500 44548
rect 24668 44380 24724 44436
rect 24444 43596 24500 43652
rect 24556 44044 24612 44100
rect 22316 40684 22372 40740
rect 22316 40348 22372 40404
rect 22428 43372 22484 43428
rect 22204 40012 22260 40068
rect 21644 39506 21700 39508
rect 21644 39454 21646 39506
rect 21646 39454 21698 39506
rect 21698 39454 21700 39506
rect 21644 39452 21700 39454
rect 21980 39506 22036 39508
rect 21980 39454 21982 39506
rect 21982 39454 22034 39506
rect 22034 39454 22036 39506
rect 21980 39452 22036 39454
rect 21868 39116 21924 39172
rect 21420 38780 21476 38836
rect 21308 38668 21364 38724
rect 21532 38668 21588 38724
rect 21532 38332 21588 38388
rect 20860 37324 20916 37380
rect 20860 36988 20916 37044
rect 20972 37100 21028 37156
rect 21756 37772 21812 37828
rect 21420 35868 21476 35924
rect 21196 35644 21252 35700
rect 22204 39452 22260 39508
rect 22876 43148 22932 43204
rect 22764 41468 22820 41524
rect 22540 40514 22596 40516
rect 22540 40462 22542 40514
rect 22542 40462 22594 40514
rect 22594 40462 22596 40514
rect 22540 40460 22596 40462
rect 22652 39004 22708 39060
rect 22764 40348 22820 40404
rect 22092 37772 22148 37828
rect 22092 36876 22148 36932
rect 22764 38668 22820 38724
rect 24220 43260 24276 43316
rect 24108 43036 24164 43092
rect 23436 42924 23492 42980
rect 23212 41580 23268 41636
rect 23212 41186 23268 41188
rect 23212 41134 23214 41186
rect 23214 41134 23266 41186
rect 23266 41134 23268 41186
rect 23212 41132 23268 41134
rect 22988 40684 23044 40740
rect 22428 38220 22484 38276
rect 23100 40460 23156 40516
rect 22988 38834 23044 38836
rect 22988 38782 22990 38834
rect 22990 38782 23042 38834
rect 23042 38782 23044 38834
rect 22988 38780 23044 38782
rect 22876 38220 22932 38276
rect 22764 38108 22820 38164
rect 22540 37490 22596 37492
rect 22540 37438 22542 37490
rect 22542 37438 22594 37490
rect 22594 37438 22596 37490
rect 22540 37436 22596 37438
rect 22988 38162 23044 38164
rect 22988 38110 22990 38162
rect 22990 38110 23042 38162
rect 23042 38110 23044 38162
rect 22988 38108 23044 38110
rect 23548 41580 23604 41636
rect 23548 40348 23604 40404
rect 24108 42364 24164 42420
rect 23996 41468 24052 41524
rect 23772 41074 23828 41076
rect 23772 41022 23774 41074
rect 23774 41022 23826 41074
rect 23826 41022 23828 41074
rect 23772 41020 23828 41022
rect 23772 40124 23828 40180
rect 24108 41020 24164 41076
rect 23996 40908 24052 40964
rect 24108 40796 24164 40852
rect 24556 42754 24612 42756
rect 24556 42702 24558 42754
rect 24558 42702 24610 42754
rect 24610 42702 24612 42754
rect 24556 42700 24612 42702
rect 24780 43650 24836 43652
rect 24780 43598 24782 43650
rect 24782 43598 24834 43650
rect 24834 43598 24836 43650
rect 24780 43596 24836 43598
rect 25340 46002 25396 46004
rect 25340 45950 25342 46002
rect 25342 45950 25394 46002
rect 25394 45950 25396 46002
rect 25340 45948 25396 45950
rect 25228 45836 25284 45892
rect 24892 42924 24948 42980
rect 25004 44380 25060 44436
rect 25340 44716 25396 44772
rect 25116 43708 25172 43764
rect 25004 43260 25060 43316
rect 25004 42700 25060 42756
rect 25116 43036 25172 43092
rect 25004 42530 25060 42532
rect 25004 42478 25006 42530
rect 25006 42478 25058 42530
rect 25058 42478 25060 42530
rect 25004 42476 25060 42478
rect 24780 41858 24836 41860
rect 24780 41806 24782 41858
rect 24782 41806 24834 41858
rect 24834 41806 24836 41858
rect 24780 41804 24836 41806
rect 24668 41468 24724 41524
rect 24780 41356 24836 41412
rect 25004 41468 25060 41524
rect 24332 40796 24388 40852
rect 24668 40684 24724 40740
rect 23996 40348 24052 40404
rect 23996 39618 24052 39620
rect 23996 39566 23998 39618
rect 23998 39566 24050 39618
rect 24050 39566 24052 39618
rect 23996 39564 24052 39566
rect 24332 39340 24388 39396
rect 24332 39058 24388 39060
rect 24332 39006 24334 39058
rect 24334 39006 24386 39058
rect 24386 39006 24388 39058
rect 24332 39004 24388 39006
rect 23436 38050 23492 38052
rect 23436 37998 23438 38050
rect 23438 37998 23490 38050
rect 23490 37998 23492 38050
rect 23436 37996 23492 37998
rect 23212 37884 23268 37940
rect 22988 37490 23044 37492
rect 22988 37438 22990 37490
rect 22990 37438 23042 37490
rect 23042 37438 23044 37490
rect 22988 37436 23044 37438
rect 23772 36764 23828 36820
rect 24780 37660 24836 37716
rect 24892 40012 24948 40068
rect 25116 39564 25172 39620
rect 25676 46284 25732 46340
rect 25452 43036 25508 43092
rect 25900 45724 25956 45780
rect 25564 42812 25620 42868
rect 25564 42642 25620 42644
rect 25564 42590 25566 42642
rect 25566 42590 25618 42642
rect 25618 42590 25620 42642
rect 25564 42588 25620 42590
rect 25452 42476 25508 42532
rect 25228 41468 25284 41524
rect 24892 37436 24948 37492
rect 25340 41804 25396 41860
rect 25340 40796 25396 40852
rect 25340 40012 25396 40068
rect 25564 42364 25620 42420
rect 25676 42028 25732 42084
rect 29372 47964 29428 48020
rect 26908 45724 26964 45780
rect 27020 47852 27076 47908
rect 26236 45612 26292 45668
rect 27356 47516 27412 47572
rect 27244 47292 27300 47348
rect 27132 46172 27188 46228
rect 27132 45500 27188 45556
rect 26124 45106 26180 45108
rect 26124 45054 26126 45106
rect 26126 45054 26178 45106
rect 26178 45054 26180 45106
rect 26124 45052 26180 45054
rect 26012 44716 26068 44772
rect 26236 44210 26292 44212
rect 26236 44158 26238 44210
rect 26238 44158 26290 44210
rect 26290 44158 26292 44210
rect 26236 44156 26292 44158
rect 26012 44044 26068 44100
rect 26012 43260 26068 43316
rect 25676 41244 25732 41300
rect 25340 39788 25396 39844
rect 26684 44828 26740 44884
rect 26796 44322 26852 44324
rect 26796 44270 26798 44322
rect 26798 44270 26850 44322
rect 26850 44270 26852 44322
rect 26796 44268 26852 44270
rect 29036 47404 29092 47460
rect 28364 47180 28420 47236
rect 27468 46732 27524 46788
rect 27468 46060 27524 46116
rect 28252 46508 28308 46564
rect 28252 45890 28308 45892
rect 28252 45838 28254 45890
rect 28254 45838 28306 45890
rect 28306 45838 28308 45890
rect 28252 45836 28308 45838
rect 27356 45218 27412 45220
rect 27356 45166 27358 45218
rect 27358 45166 27410 45218
rect 27410 45166 27412 45218
rect 27356 45164 27412 45166
rect 27692 44828 27748 44884
rect 27692 44380 27748 44436
rect 27356 44322 27412 44324
rect 27356 44270 27358 44322
rect 27358 44270 27410 44322
rect 27410 44270 27412 44322
rect 27356 44268 27412 44270
rect 26348 43372 26404 43428
rect 26684 44044 26740 44100
rect 26236 42700 26292 42756
rect 26124 42530 26180 42532
rect 26124 42478 26126 42530
rect 26126 42478 26178 42530
rect 26178 42478 26180 42530
rect 26124 42476 26180 42478
rect 26236 41186 26292 41188
rect 26236 41134 26238 41186
rect 26238 41134 26290 41186
rect 26290 41134 26292 41186
rect 26236 41132 26292 41134
rect 26012 40402 26068 40404
rect 26012 40350 26014 40402
rect 26014 40350 26066 40402
rect 26066 40350 26068 40402
rect 26012 40348 26068 40350
rect 26460 41692 26516 41748
rect 26460 40796 26516 40852
rect 26348 40124 26404 40180
rect 25788 39618 25844 39620
rect 25788 39566 25790 39618
rect 25790 39566 25842 39618
rect 25842 39566 25844 39618
rect 25788 39564 25844 39566
rect 25452 39452 25508 39508
rect 25228 36428 25284 36484
rect 24668 36316 24724 36372
rect 22540 35532 22596 35588
rect 27692 43708 27748 43764
rect 26796 43484 26852 43540
rect 27244 43484 27300 43540
rect 26684 42588 26740 42644
rect 27020 42978 27076 42980
rect 27020 42926 27022 42978
rect 27022 42926 27074 42978
rect 27074 42926 27076 42978
rect 27020 42924 27076 42926
rect 27132 42866 27188 42868
rect 27132 42814 27134 42866
rect 27134 42814 27186 42866
rect 27186 42814 27188 42866
rect 27132 42812 27188 42814
rect 26796 42476 26852 42532
rect 26684 41692 26740 41748
rect 26572 36988 26628 37044
rect 27020 42588 27076 42644
rect 26908 42364 26964 42420
rect 27916 43596 27972 43652
rect 27804 43538 27860 43540
rect 27804 43486 27806 43538
rect 27806 43486 27858 43538
rect 27858 43486 27860 43538
rect 27804 43484 27860 43486
rect 27580 42866 27636 42868
rect 27580 42814 27582 42866
rect 27582 42814 27634 42866
rect 27634 42814 27636 42866
rect 27580 42812 27636 42814
rect 27468 42700 27524 42756
rect 27020 38780 27076 38836
rect 27356 40626 27412 40628
rect 27356 40574 27358 40626
rect 27358 40574 27410 40626
rect 27410 40574 27412 40626
rect 27356 40572 27412 40574
rect 27020 38332 27076 38388
rect 27916 43148 27972 43204
rect 28364 44940 28420 44996
rect 28140 44604 28196 44660
rect 28364 44604 28420 44660
rect 28140 44044 28196 44100
rect 28028 42812 28084 42868
rect 28140 43820 28196 43876
rect 28028 42530 28084 42532
rect 28028 42478 28030 42530
rect 28030 42478 28082 42530
rect 28082 42478 28084 42530
rect 28028 42476 28084 42478
rect 27692 42140 27748 42196
rect 28028 41468 28084 41524
rect 28924 44604 28980 44660
rect 28588 44098 28644 44100
rect 28588 44046 28590 44098
rect 28590 44046 28642 44098
rect 28642 44046 28644 44098
rect 28588 44044 28644 44046
rect 28588 43820 28644 43876
rect 28924 43708 28980 43764
rect 30044 47740 30100 47796
rect 29372 45052 29428 45108
rect 29372 44492 29428 44548
rect 29596 45666 29652 45668
rect 29596 45614 29598 45666
rect 29598 45614 29650 45666
rect 29650 45614 29652 45666
rect 29596 45612 29652 45614
rect 29484 44380 29540 44436
rect 29596 44940 29652 44996
rect 29148 43820 29204 43876
rect 28364 43260 28420 43316
rect 29372 43538 29428 43540
rect 29372 43486 29374 43538
rect 29374 43486 29426 43538
rect 29426 43486 29428 43538
rect 29372 43484 29428 43486
rect 29148 43148 29204 43204
rect 28476 43036 28532 43092
rect 28252 42252 28308 42308
rect 29484 42252 29540 42308
rect 33180 47068 33236 47124
rect 32284 45948 32340 46004
rect 32396 46060 32452 46116
rect 30380 45778 30436 45780
rect 30380 45726 30382 45778
rect 30382 45726 30434 45778
rect 30434 45726 30436 45778
rect 30380 45724 30436 45726
rect 30604 45500 30660 45556
rect 29932 44994 29988 44996
rect 29932 44942 29934 44994
rect 29934 44942 29986 44994
rect 29986 44942 29988 44994
rect 29932 44940 29988 44942
rect 29932 44322 29988 44324
rect 29932 44270 29934 44322
rect 29934 44270 29986 44322
rect 29986 44270 29988 44322
rect 29932 44268 29988 44270
rect 29820 44156 29876 44212
rect 30044 44156 30100 44212
rect 29820 43260 29876 43316
rect 30716 45388 30772 45444
rect 30828 44604 30884 44660
rect 30380 44210 30436 44212
rect 30380 44158 30382 44210
rect 30382 44158 30434 44210
rect 30434 44158 30436 44210
rect 30380 44156 30436 44158
rect 30716 44044 30772 44100
rect 30268 43148 30324 43204
rect 29596 42140 29652 42196
rect 28476 41468 28532 41524
rect 31052 45500 31108 45556
rect 31948 45890 32004 45892
rect 31948 45838 31950 45890
rect 31950 45838 32002 45890
rect 32002 45838 32004 45890
rect 31948 45836 32004 45838
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 33852 46002 33908 46004
rect 33852 45950 33854 46002
rect 33854 45950 33906 46002
rect 33906 45950 33908 46002
rect 33852 45948 33908 45950
rect 31724 45388 31780 45444
rect 31612 45218 31668 45220
rect 31612 45166 31614 45218
rect 31614 45166 31666 45218
rect 31666 45166 31668 45218
rect 31612 45164 31668 45166
rect 34748 45330 34804 45332
rect 34748 45278 34750 45330
rect 34750 45278 34802 45330
rect 34802 45278 34804 45330
rect 34748 45276 34804 45278
rect 42476 46396 42532 46452
rect 43036 45948 43092 46004
rect 43708 46002 43764 46004
rect 43708 45950 43710 46002
rect 43710 45950 43762 46002
rect 43762 45950 43764 46002
rect 43708 45948 43764 45950
rect 35084 45276 35140 45332
rect 32508 45106 32564 45108
rect 32508 45054 32510 45106
rect 32510 45054 32562 45106
rect 32562 45054 32564 45106
rect 32508 45052 32564 45054
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 32172 44434 32228 44436
rect 32172 44382 32174 44434
rect 32174 44382 32226 44434
rect 32226 44382 32228 44434
rect 32172 44380 32228 44382
rect 32060 43596 32116 43652
rect 31276 43372 31332 43428
rect 30940 41804 30996 41860
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 32620 40572 32676 40628
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 48076 39676 48132 39732
rect 29372 38892 29428 38948
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 48076 37660 48132 37716
rect 27916 36764 27972 36820
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 27468 36540 27524 36596
rect 26796 35756 26852 35812
rect 48076 35644 48132 35700
rect 26236 35196 26292 35252
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 21868 34972 21924 35028
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 48076 34300 48132 34356
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 19628 33516 19684 33572
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 48076 32284 48132 32340
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 48076 30940 48132 30996
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 48076 28924 48132 28980
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 48076 26850 48132 26852
rect 48076 26798 48078 26850
rect 48078 26798 48130 26850
rect 48130 26798 48132 26850
rect 48076 26796 48132 26798
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 48076 23548 48132 23604
rect 20044 23492 20100 23494
rect 11228 23324 11284 23380
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 48076 21532 48132 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 48076 18562 48132 18564
rect 48076 18510 48078 18562
rect 48078 18510 48130 18562
rect 48130 18510 48132 18562
rect 48076 18508 48132 18510
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 48076 16828 48132 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 48076 12850 48132 12852
rect 48076 12798 48078 12850
rect 48078 12798 48130 12850
rect 48130 12798 48132 12850
rect 48076 12796 48132 12798
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 48076 11452 48132 11508
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 48076 9436 48132 9492
rect 20044 9380 20100 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 48076 7420 48132 7476
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 48076 6076 48132 6132
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 5852 3612 5908 3668
rect 2492 2268 2548 2324
rect 4732 3276 4788 3332
rect 5740 3330 5796 3332
rect 5740 3278 5742 3330
rect 5742 3278 5794 3330
rect 5794 3278 5796 3330
rect 5740 3276 5796 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 28252 3276 28308 3332
rect 29260 3330 29316 3332
rect 29260 3278 29262 3330
rect 29262 3278 29314 3330
rect 29314 3278 29316 3330
rect 29260 3276 29316 3278
rect 47404 2044 47460 2100
rect 48076 700 48132 756
<< metal3 >>
rect 200 49140 800 49168
rect 200 49084 3388 49140
rect 3444 49084 3454 49140
rect 200 49056 800 49084
rect 49200 48384 49800 48496
rect 11330 48188 11340 48244
rect 11396 48188 24220 48244
rect 24276 48188 24286 48244
rect 10658 48076 10668 48132
rect 10724 48076 25452 48132
rect 25508 48076 25518 48132
rect 16706 47964 16716 48020
rect 16772 47964 29372 48020
rect 29428 47964 29438 48020
rect 14018 47852 14028 47908
rect 14084 47852 27020 47908
rect 27076 47852 27086 47908
rect 200 47712 800 47824
rect 9986 47740 9996 47796
rect 10052 47740 30044 47796
rect 30100 47740 30110 47796
rect 10882 47628 10892 47684
rect 10948 47628 11452 47684
rect 11508 47628 11518 47684
rect 15698 47516 15708 47572
rect 15764 47516 27356 47572
rect 27412 47516 27422 47572
rect 16594 47404 16604 47460
rect 16660 47404 29036 47460
rect 29092 47404 29102 47460
rect 16034 47292 16044 47348
rect 16100 47292 27244 47348
rect 27300 47292 27310 47348
rect 20290 47180 20300 47236
rect 20356 47180 28364 47236
rect 28420 47180 28430 47236
rect 20514 47068 20524 47124
rect 20580 47068 33180 47124
rect 33236 47068 33246 47124
rect 19394 46732 19404 46788
rect 19460 46732 27468 46788
rect 27524 46732 27534 46788
rect 12786 46508 12796 46564
rect 12852 46508 24892 46564
rect 24948 46508 28252 46564
rect 28308 46508 28318 46564
rect 3042 46396 3052 46452
rect 3108 46396 12236 46452
rect 12292 46396 12302 46452
rect 24434 46396 24444 46452
rect 24500 46396 42476 46452
rect 42532 46396 42542 46452
rect 49200 46368 49800 46480
rect 14130 46284 14140 46340
rect 14196 46284 25676 46340
rect 25732 46284 25742 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 16258 46172 16268 46228
rect 16324 46172 27132 46228
rect 27188 46172 27198 46228
rect 6850 46060 6860 46116
rect 6916 46060 24668 46116
rect 24724 46060 24734 46116
rect 27458 46060 27468 46116
rect 27524 46060 32396 46116
rect 32452 46060 32462 46116
rect 7970 45948 7980 46004
rect 8036 45948 12572 46004
rect 12628 45948 12638 46004
rect 17612 45948 20300 46004
rect 20356 45948 20366 46004
rect 21074 45948 21084 46004
rect 21140 45948 25340 46004
rect 25396 45948 25406 46004
rect 32274 45948 32284 46004
rect 32340 45948 33852 46004
rect 33908 45948 33918 46004
rect 43026 45948 43036 46004
rect 43092 45948 43708 46004
rect 43764 45948 43774 46004
rect 4946 45836 4956 45892
rect 5012 45836 13580 45892
rect 13636 45836 13646 45892
rect 14466 45836 14476 45892
rect 14532 45836 15932 45892
rect 15988 45836 15998 45892
rect 200 45780 800 45808
rect 17612 45780 17668 45948
rect 19954 45836 19964 45892
rect 20020 45836 25228 45892
rect 25284 45836 25294 45892
rect 28242 45836 28252 45892
rect 28308 45836 31948 45892
rect 32004 45836 32014 45892
rect 200 45724 2492 45780
rect 2548 45724 2558 45780
rect 8054 45724 8092 45780
rect 8148 45724 8158 45780
rect 9538 45724 9548 45780
rect 9604 45724 10892 45780
rect 10948 45724 10958 45780
rect 12114 45724 12124 45780
rect 12180 45724 17668 45780
rect 17826 45724 17836 45780
rect 17892 45724 25900 45780
rect 25956 45724 25966 45780
rect 26898 45724 26908 45780
rect 26964 45724 30380 45780
rect 30436 45724 30446 45780
rect 200 45696 800 45724
rect 1810 45612 1820 45668
rect 1876 45612 3500 45668
rect 3556 45612 4284 45668
rect 4340 45612 4350 45668
rect 5506 45612 5516 45668
rect 5572 45612 16380 45668
rect 16436 45612 16446 45668
rect 17490 45612 17500 45668
rect 17556 45612 18956 45668
rect 19012 45612 19022 45668
rect 26226 45612 26236 45668
rect 26292 45612 29596 45668
rect 29652 45612 29662 45668
rect 4162 45500 4172 45556
rect 4228 45500 10668 45556
rect 10724 45500 10734 45556
rect 10994 45500 11004 45556
rect 11060 45500 12404 45556
rect 12562 45500 12572 45556
rect 12628 45500 19628 45556
rect 19684 45500 19694 45556
rect 22082 45500 22092 45556
rect 22148 45500 24444 45556
rect 24500 45500 24510 45556
rect 27122 45500 27132 45556
rect 27188 45500 30604 45556
rect 30660 45500 31052 45556
rect 31108 45500 31118 45556
rect 12348 45444 12404 45500
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 5730 45388 5740 45444
rect 5796 45388 12124 45444
rect 12180 45388 12190 45444
rect 12348 45388 18396 45444
rect 18452 45388 18462 45444
rect 24210 45388 24220 45444
rect 24276 45388 30716 45444
rect 30772 45388 31724 45444
rect 31780 45388 31790 45444
rect 3154 45276 3164 45332
rect 3220 45276 9996 45332
rect 10052 45276 10062 45332
rect 14914 45276 14924 45332
rect 14980 45276 15372 45332
rect 15428 45276 16492 45332
rect 16548 45276 20636 45332
rect 20692 45276 20702 45332
rect 23762 45276 23772 45332
rect 23828 45276 34748 45332
rect 34804 45276 35084 45332
rect 35140 45276 35150 45332
rect 7746 45164 7756 45220
rect 7812 45164 8988 45220
rect 9044 45164 15820 45220
rect 15876 45164 16716 45220
rect 16772 45164 16782 45220
rect 18386 45164 18396 45220
rect 18452 45164 20972 45220
rect 21028 45164 21038 45220
rect 27346 45164 27356 45220
rect 27412 45164 31612 45220
rect 31668 45164 31678 45220
rect 4274 45052 4284 45108
rect 4340 45052 6188 45108
rect 6244 45052 8764 45108
rect 8820 45052 8830 45108
rect 10070 45052 10108 45108
rect 10164 45052 10174 45108
rect 11106 45052 11116 45108
rect 11172 45052 14588 45108
rect 14644 45052 14654 45108
rect 16342 45052 16380 45108
rect 16436 45052 16446 45108
rect 21410 45052 21420 45108
rect 21476 45052 26124 45108
rect 26180 45052 26190 45108
rect 29362 45052 29372 45108
rect 29428 45052 32508 45108
rect 32564 45052 32574 45108
rect 49200 45024 49800 45136
rect 4946 44940 4956 44996
rect 5012 44940 9548 44996
rect 9604 44940 9614 44996
rect 11442 44940 11452 44996
rect 11508 44940 15932 44996
rect 15988 44940 15998 44996
rect 28354 44940 28364 44996
rect 28420 44940 29596 44996
rect 29652 44940 29932 44996
rect 29988 44940 29998 44996
rect 9650 44828 9660 44884
rect 9716 44828 11676 44884
rect 11732 44828 14588 44884
rect 14644 44828 14654 44884
rect 26674 44828 26684 44884
rect 26740 44828 27692 44884
rect 27748 44828 27758 44884
rect 10994 44716 11004 44772
rect 11060 44716 16492 44772
rect 16548 44716 16558 44772
rect 20850 44716 20860 44772
rect 20916 44716 21308 44772
rect 21364 44716 22540 44772
rect 22596 44716 22606 44772
rect 25330 44716 25340 44772
rect 25396 44716 26012 44772
rect 26068 44716 26078 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 8866 44604 8876 44660
rect 8932 44604 21756 44660
rect 21812 44604 21822 44660
rect 22306 44604 22316 44660
rect 22372 44604 28140 44660
rect 28196 44604 28206 44660
rect 28354 44604 28364 44660
rect 28420 44604 28924 44660
rect 28980 44604 30828 44660
rect 30884 44604 30894 44660
rect 7858 44492 7868 44548
rect 7924 44492 11228 44548
rect 11284 44492 11564 44548
rect 11620 44492 11630 44548
rect 19618 44492 19628 44548
rect 19684 44492 24444 44548
rect 24500 44492 24510 44548
rect 27132 44492 29372 44548
rect 29428 44492 29438 44548
rect 3714 44380 3724 44436
rect 3780 44380 11004 44436
rect 11060 44380 11070 44436
rect 15138 44380 15148 44436
rect 15204 44380 15596 44436
rect 15652 44380 22428 44436
rect 22484 44380 22494 44436
rect 24658 44380 24668 44436
rect 24724 44380 25004 44436
rect 25060 44380 25070 44436
rect 5842 44268 5852 44324
rect 5908 44268 6524 44324
rect 6580 44268 6590 44324
rect 10434 44268 10444 44324
rect 10500 44268 16828 44324
rect 16884 44268 16894 44324
rect 17042 44268 17052 44324
rect 17108 44268 26796 44324
rect 26852 44268 26862 44324
rect 27132 44212 27188 44492
rect 27682 44380 27692 44436
rect 27748 44380 29484 44436
rect 29540 44380 32172 44436
rect 32228 44380 32238 44436
rect 27346 44268 27356 44324
rect 27412 44268 29932 44324
rect 29988 44268 29998 44324
rect 7298 44156 7308 44212
rect 7364 44156 11228 44212
rect 11284 44156 11294 44212
rect 11442 44156 11452 44212
rect 11508 44156 15820 44212
rect 15876 44156 16156 44212
rect 16212 44156 16222 44212
rect 17378 44156 17388 44212
rect 17444 44156 20860 44212
rect 20916 44156 20926 44212
rect 26226 44156 26236 44212
rect 26292 44156 27188 44212
rect 27916 44156 29820 44212
rect 29876 44156 30044 44212
rect 30100 44156 30380 44212
rect 30436 44156 30446 44212
rect 27916 44100 27972 44156
rect 4610 44044 4620 44100
rect 4676 44044 14140 44100
rect 14196 44044 15148 44100
rect 16258 44044 16268 44100
rect 16324 44044 20188 44100
rect 20244 44044 20254 44100
rect 20626 44044 20636 44100
rect 20692 44044 24556 44100
rect 24612 44044 24622 44100
rect 26002 44044 26012 44100
rect 26068 44044 26684 44100
rect 26740 44044 26750 44100
rect 26898 44044 26908 44100
rect 26964 44044 27972 44100
rect 28130 44044 28140 44100
rect 28196 44044 28588 44100
rect 28644 44044 30716 44100
rect 30772 44044 30782 44100
rect 15092 43988 15148 44044
rect 5058 43932 5068 43988
rect 5124 43932 10668 43988
rect 10724 43932 11452 43988
rect 11508 43932 11518 43988
rect 15092 43932 18172 43988
rect 18228 43932 19180 43988
rect 19236 43932 19246 43988
rect 22418 43932 22428 43988
rect 22484 43932 28420 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 4050 43820 4060 43876
rect 4116 43820 5180 43876
rect 5236 43820 5246 43876
rect 6738 43820 6748 43876
rect 6804 43820 7420 43876
rect 7476 43820 7486 43876
rect 20626 43820 20636 43876
rect 20692 43820 26740 43876
rect 26796 43820 26908 43932
rect 28364 43876 28420 43932
rect 27468 43820 28140 43876
rect 28196 43820 28206 43876
rect 28364 43820 28588 43876
rect 28644 43820 29148 43876
rect 29204 43820 29214 43876
rect 200 43764 800 43792
rect 20636 43764 20692 43820
rect 26684 43764 26740 43820
rect 27468 43764 27524 43820
rect 200 43708 2156 43764
rect 2212 43708 2222 43764
rect 4834 43708 4844 43764
rect 4900 43708 7868 43764
rect 7924 43708 7934 43764
rect 8978 43708 8988 43764
rect 9044 43708 9660 43764
rect 9716 43708 9726 43764
rect 10098 43708 10108 43764
rect 10164 43708 10332 43764
rect 10388 43708 10398 43764
rect 16818 43708 16828 43764
rect 16884 43708 20692 43764
rect 21634 43708 21644 43764
rect 21700 43708 25116 43764
rect 25172 43708 25182 43764
rect 26684 43708 27524 43764
rect 27682 43708 27692 43764
rect 27748 43708 28924 43764
rect 28980 43708 28990 43764
rect 200 43680 800 43708
rect 5058 43596 5068 43652
rect 5124 43596 6076 43652
rect 6132 43596 8876 43652
rect 8932 43596 9100 43652
rect 9156 43596 9166 43652
rect 16930 43596 16940 43652
rect 16996 43596 24276 43652
rect 24434 43596 24444 43652
rect 24500 43596 24780 43652
rect 24836 43596 24846 43652
rect 27906 43596 27916 43652
rect 27972 43596 32060 43652
rect 32116 43596 32126 43652
rect 24220 43540 24276 43596
rect 5170 43484 5180 43540
rect 5236 43484 8764 43540
rect 8820 43484 13692 43540
rect 13748 43484 13758 43540
rect 14018 43484 14028 43540
rect 14084 43484 21644 43540
rect 21700 43484 21980 43540
rect 22036 43484 22046 43540
rect 24220 43484 25284 43540
rect 26786 43484 26796 43540
rect 26852 43484 26862 43540
rect 27234 43484 27244 43540
rect 27300 43484 27804 43540
rect 27860 43484 29372 43540
rect 29428 43484 29438 43540
rect 25228 43428 25284 43484
rect 26796 43428 26852 43484
rect 3490 43372 3500 43428
rect 3556 43372 5404 43428
rect 5460 43372 5470 43428
rect 7298 43372 7308 43428
rect 7364 43372 8540 43428
rect 8596 43372 8606 43428
rect 8838 43372 8876 43428
rect 8932 43372 8942 43428
rect 12562 43372 12572 43428
rect 12628 43372 13468 43428
rect 13524 43372 13534 43428
rect 19618 43372 19628 43428
rect 19684 43372 21196 43428
rect 21252 43372 21262 43428
rect 21522 43372 21532 43428
rect 21588 43372 22428 43428
rect 22484 43372 22494 43428
rect 25228 43372 26348 43428
rect 26404 43372 31276 43428
rect 31332 43372 31342 43428
rect 15698 43260 15708 43316
rect 15764 43260 16604 43316
rect 16660 43260 16670 43316
rect 16818 43260 16828 43316
rect 16884 43260 24220 43316
rect 24276 43260 24286 43316
rect 24994 43260 25004 43316
rect 25060 43260 26012 43316
rect 26068 43260 28364 43316
rect 28420 43260 29820 43316
rect 29876 43260 29886 43316
rect 13682 43148 13692 43204
rect 13748 43148 17724 43204
rect 17780 43148 18172 43204
rect 18228 43148 18238 43204
rect 22866 43148 22876 43204
rect 22932 43148 27916 43204
rect 27972 43148 27982 43204
rect 29138 43148 29148 43204
rect 29204 43148 30268 43204
rect 30324 43148 30334 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 8418 43036 8428 43092
rect 8484 43036 9324 43092
rect 9380 43036 10556 43092
rect 10612 43036 14364 43092
rect 14420 43036 15708 43092
rect 15764 43036 15774 43092
rect 16146 43036 16156 43092
rect 16212 43036 21868 43092
rect 21924 43036 21934 43092
rect 24098 43036 24108 43092
rect 24164 43036 25116 43092
rect 25172 43036 25182 43092
rect 25442 43036 25452 43092
rect 25508 43036 26628 43092
rect 26786 43036 26796 43092
rect 26852 43036 28476 43092
rect 28532 43036 28542 43092
rect 26572 42980 26628 43036
rect 49200 43008 49800 43120
rect 6626 42924 6636 42980
rect 6692 42924 11340 42980
rect 11396 42924 11406 42980
rect 11554 42924 11564 42980
rect 11620 42924 13916 42980
rect 13972 42924 13982 42980
rect 15250 42924 15260 42980
rect 15316 42924 20860 42980
rect 20916 42924 20926 42980
rect 21186 42924 21196 42980
rect 21252 42924 23436 42980
rect 23492 42924 23502 42980
rect 24882 42924 24892 42980
rect 24948 42924 26516 42980
rect 26572 42924 27020 42980
rect 27076 42924 27086 42980
rect 26460 42868 26516 42924
rect 3938 42812 3948 42868
rect 4004 42812 4508 42868
rect 4564 42812 7308 42868
rect 7364 42812 7374 42868
rect 7634 42812 7644 42868
rect 7700 42812 7980 42868
rect 8036 42812 8046 42868
rect 10210 42812 10220 42868
rect 10276 42812 15708 42868
rect 15764 42812 15774 42868
rect 16034 42812 16044 42868
rect 16100 42812 18620 42868
rect 18676 42812 20076 42868
rect 20132 42812 20468 42868
rect 20738 42812 20748 42868
rect 20804 42812 25564 42868
rect 25620 42812 25630 42868
rect 26460 42812 27132 42868
rect 27188 42812 27580 42868
rect 27636 42812 27646 42868
rect 28018 42812 28028 42868
rect 28084 42812 28094 42868
rect 7074 42700 7084 42756
rect 7140 42700 8204 42756
rect 8260 42700 8270 42756
rect 9426 42700 9436 42756
rect 9492 42700 9884 42756
rect 9940 42700 9950 42756
rect 10098 42700 10108 42756
rect 10164 42700 14364 42756
rect 14420 42700 14430 42756
rect 14364 42644 14420 42700
rect 20412 42644 20468 42812
rect 28028 42756 28084 42812
rect 24546 42700 24556 42756
rect 24612 42700 25004 42756
rect 25060 42700 25070 42756
rect 25228 42700 25844 42756
rect 26226 42700 26236 42756
rect 26292 42700 26796 42756
rect 26852 42700 26862 42756
rect 27458 42700 27468 42756
rect 27524 42700 28084 42756
rect 25228 42644 25284 42700
rect 25788 42644 25844 42700
rect 8306 42588 8316 42644
rect 8372 42588 8652 42644
rect 8708 42588 9996 42644
rect 10052 42588 10062 42644
rect 14364 42588 15036 42644
rect 15092 42588 15102 42644
rect 20412 42588 25284 42644
rect 25526 42588 25564 42644
rect 25620 42588 25630 42644
rect 25788 42588 26404 42644
rect 26674 42588 26684 42644
rect 26740 42588 27020 42644
rect 27076 42588 27086 42644
rect 8082 42476 8092 42532
rect 8148 42476 10780 42532
rect 10836 42476 10846 42532
rect 11442 42476 11452 42532
rect 11508 42476 12908 42532
rect 12964 42476 14924 42532
rect 14980 42476 14990 42532
rect 16594 42476 16604 42532
rect 16660 42476 20244 42532
rect 20822 42476 20860 42532
rect 20916 42476 20926 42532
rect 24966 42476 25004 42532
rect 25060 42476 25070 42532
rect 25442 42476 25452 42532
rect 25508 42476 26124 42532
rect 26180 42476 26190 42532
rect 200 42420 800 42448
rect 20188 42420 20244 42476
rect 26348 42420 26404 42588
rect 26786 42476 26796 42532
rect 26852 42476 28028 42532
rect 28084 42476 28094 42532
rect 200 42364 1820 42420
rect 1876 42364 1886 42420
rect 9986 42364 9996 42420
rect 10052 42364 11564 42420
rect 11620 42364 12124 42420
rect 12180 42364 12190 42420
rect 13906 42364 13916 42420
rect 13972 42364 16044 42420
rect 16100 42364 16110 42420
rect 20188 42364 21980 42420
rect 22036 42364 24108 42420
rect 24164 42364 25564 42420
rect 25620 42364 25630 42420
rect 26348 42364 26908 42420
rect 26964 42364 26974 42420
rect 200 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 13794 42252 13804 42308
rect 13860 42252 18060 42308
rect 18116 42252 18126 42308
rect 20290 42252 20300 42308
rect 20356 42252 28252 42308
rect 28308 42252 29484 42308
rect 29540 42252 29550 42308
rect 4274 42140 4284 42196
rect 4340 42140 5628 42196
rect 5684 42140 5694 42196
rect 6178 42140 6188 42196
rect 6244 42140 8316 42196
rect 8372 42140 8382 42196
rect 8754 42140 8764 42196
rect 8820 42140 10892 42196
rect 10948 42140 10958 42196
rect 14354 42140 14364 42196
rect 14420 42140 15484 42196
rect 15540 42140 15550 42196
rect 20514 42140 20524 42196
rect 20580 42140 21756 42196
rect 21812 42140 21822 42196
rect 27682 42140 27692 42196
rect 27748 42140 29596 42196
rect 29652 42140 29662 42196
rect 7522 42028 7532 42084
rect 7588 42028 11340 42084
rect 11396 42028 11406 42084
rect 12562 42028 12572 42084
rect 12628 42028 16268 42084
rect 16324 42028 16334 42084
rect 16818 42028 16828 42084
rect 16884 42028 17724 42084
rect 17780 42028 17790 42084
rect 18274 42028 18284 42084
rect 18340 42028 19964 42084
rect 20020 42028 20030 42084
rect 20626 42028 20636 42084
rect 20692 42028 25676 42084
rect 25732 42028 25742 42084
rect 6290 41916 6300 41972
rect 6356 41916 10220 41972
rect 10276 41916 18508 41972
rect 18564 41916 18574 41972
rect 7074 41804 7084 41860
rect 7140 41804 9996 41860
rect 10052 41804 10062 41860
rect 14550 41804 14588 41860
rect 14644 41804 14654 41860
rect 15810 41804 15820 41860
rect 15876 41804 16380 41860
rect 16436 41804 17052 41860
rect 17108 41804 17948 41860
rect 18004 41804 18014 41860
rect 19058 41804 19068 41860
rect 19124 41804 20748 41860
rect 20804 41804 22092 41860
rect 22148 41804 22158 41860
rect 24770 41804 24780 41860
rect 24836 41804 25340 41860
rect 25396 41804 30940 41860
rect 30996 41804 31006 41860
rect 6066 41692 6076 41748
rect 6132 41692 7420 41748
rect 7476 41692 7486 41748
rect 8092 41692 9660 41748
rect 9716 41692 13692 41748
rect 13748 41692 13758 41748
rect 14466 41692 14476 41748
rect 14532 41692 18060 41748
rect 18116 41692 18126 41748
rect 26450 41692 26460 41748
rect 26516 41692 26684 41748
rect 26740 41692 26750 41748
rect 8092 41636 8148 41692
rect 4946 41580 4956 41636
rect 5012 41580 8092 41636
rect 8148 41580 8158 41636
rect 8642 41580 8652 41636
rect 8708 41580 15148 41636
rect 15204 41580 15214 41636
rect 15586 41580 15596 41636
rect 15652 41580 16156 41636
rect 16212 41580 16222 41636
rect 16370 41580 16380 41636
rect 16436 41580 20300 41636
rect 20356 41580 23212 41636
rect 23268 41580 23548 41636
rect 23604 41580 23614 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 7298 41468 7308 41524
rect 7364 41468 10332 41524
rect 10388 41468 10398 41524
rect 11330 41468 11340 41524
rect 11396 41468 16604 41524
rect 16660 41468 17836 41524
rect 17892 41468 17902 41524
rect 20402 41468 20412 41524
rect 20468 41468 20860 41524
rect 20916 41468 22764 41524
rect 22820 41468 23996 41524
rect 24052 41468 24062 41524
rect 24658 41468 24668 41524
rect 24724 41468 25004 41524
rect 25060 41468 25070 41524
rect 25218 41468 25228 41524
rect 25284 41468 28028 41524
rect 28084 41468 28476 41524
rect 28532 41468 28542 41524
rect 7970 41356 7980 41412
rect 8036 41356 12908 41412
rect 12964 41356 13244 41412
rect 13300 41356 13310 41412
rect 14914 41356 14924 41412
rect 14980 41356 15018 41412
rect 15138 41356 15148 41412
rect 15204 41356 16380 41412
rect 16436 41356 16446 41412
rect 17714 41356 17724 41412
rect 17780 41356 20524 41412
rect 20580 41356 24780 41412
rect 24836 41356 24846 41412
rect 6402 41244 6412 41300
rect 6468 41244 8092 41300
rect 8148 41244 8158 41300
rect 9538 41244 9548 41300
rect 9604 41244 16716 41300
rect 16772 41244 16782 41300
rect 18722 41244 18732 41300
rect 18788 41244 25676 41300
rect 25732 41244 25742 41300
rect 9090 41132 9100 41188
rect 9156 41132 10108 41188
rect 10164 41132 11676 41188
rect 11732 41132 11742 41188
rect 13682 41132 13692 41188
rect 13748 41132 15820 41188
rect 15876 41132 15886 41188
rect 16146 41132 16156 41188
rect 16212 41132 20300 41188
rect 20356 41132 20366 41188
rect 20626 41132 20636 41188
rect 20692 41132 21196 41188
rect 21252 41132 21262 41188
rect 21746 41132 21756 41188
rect 21812 41132 22988 41188
rect 23044 41132 23212 41188
rect 23268 41132 25564 41188
rect 25620 41132 26236 41188
rect 26292 41132 26302 41188
rect 5618 41020 5628 41076
rect 5684 41020 9996 41076
rect 10052 41020 10062 41076
rect 11442 41020 11452 41076
rect 11508 41020 15484 41076
rect 15540 41020 16380 41076
rect 16436 41020 16446 41076
rect 18508 41020 19628 41076
rect 19684 41020 20748 41076
rect 20804 41020 20814 41076
rect 22082 41020 22092 41076
rect 22148 41020 23772 41076
rect 23828 41020 23838 41076
rect 24098 41020 24108 41076
rect 24164 41020 26908 41076
rect 9996 40964 10052 41020
rect 18508 40964 18564 41020
rect 9996 40908 11340 40964
rect 11396 40908 11406 40964
rect 14102 40908 14140 40964
rect 14196 40908 14206 40964
rect 14914 40908 14924 40964
rect 14980 40908 18564 40964
rect 19842 40908 19852 40964
rect 19908 40908 23996 40964
rect 24052 40908 24062 40964
rect 14802 40796 14812 40852
rect 14868 40796 17052 40852
rect 17108 40796 17118 40852
rect 21606 40796 21644 40852
rect 21700 40796 21710 40852
rect 22530 40796 22540 40852
rect 22596 40796 24108 40852
rect 24164 40796 24174 40852
rect 24322 40796 24332 40852
rect 24388 40796 25340 40852
rect 25396 40796 26460 40852
rect 26516 40796 26526 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 15810 40684 15820 40740
rect 15876 40684 16268 40740
rect 16324 40684 16334 40740
rect 16930 40684 16940 40740
rect 16996 40684 19404 40740
rect 19460 40684 19470 40740
rect 20290 40684 20300 40740
rect 20356 40684 22316 40740
rect 22372 40684 22382 40740
rect 22866 40684 22876 40740
rect 22932 40684 22988 40740
rect 23044 40684 23054 40740
rect 24658 40684 24668 40740
rect 24724 40684 24734 40740
rect 24668 40628 24724 40684
rect 9650 40572 9660 40628
rect 9716 40572 10220 40628
rect 10276 40572 14364 40628
rect 14420 40572 14430 40628
rect 15698 40572 15708 40628
rect 15764 40572 16604 40628
rect 16660 40572 16670 40628
rect 19842 40572 19852 40628
rect 19908 40572 24724 40628
rect 26852 40628 26908 41020
rect 49200 40992 49800 41104
rect 26852 40572 27356 40628
rect 27412 40572 32620 40628
rect 32676 40572 32686 40628
rect 9202 40460 9212 40516
rect 9268 40460 11340 40516
rect 11396 40460 11406 40516
rect 13682 40460 13692 40516
rect 13748 40460 16940 40516
rect 16996 40460 17006 40516
rect 19180 40460 22540 40516
rect 22596 40460 23100 40516
rect 23156 40460 23166 40516
rect 200 40320 800 40432
rect 19180 40404 19236 40460
rect 8194 40348 8204 40404
rect 8260 40348 10108 40404
rect 10164 40348 10556 40404
rect 10612 40348 10622 40404
rect 12114 40348 12124 40404
rect 12180 40348 14924 40404
rect 14980 40348 14990 40404
rect 18162 40348 18172 40404
rect 18228 40348 19180 40404
rect 19236 40348 19246 40404
rect 20402 40348 20412 40404
rect 20468 40348 20748 40404
rect 20804 40348 20814 40404
rect 20962 40348 20972 40404
rect 21028 40348 21066 40404
rect 22306 40348 22316 40404
rect 22372 40348 22764 40404
rect 22820 40348 22830 40404
rect 23538 40348 23548 40404
rect 23604 40348 23996 40404
rect 24052 40348 26012 40404
rect 26068 40348 26078 40404
rect 14354 40236 14364 40292
rect 14420 40236 17948 40292
rect 18004 40236 18014 40292
rect 20402 40236 20412 40292
rect 20468 40236 26684 40292
rect 26740 40236 26750 40292
rect 6626 40124 6636 40180
rect 6692 40124 13020 40180
rect 13076 40124 15372 40180
rect 15428 40124 15820 40180
rect 15876 40124 15886 40180
rect 18946 40124 18956 40180
rect 19012 40124 21756 40180
rect 21812 40124 23772 40180
rect 23828 40124 26348 40180
rect 26404 40124 26414 40180
rect 8306 40012 8316 40068
rect 8372 40012 12348 40068
rect 12404 40012 15596 40068
rect 15652 40012 15662 40068
rect 16370 40012 16380 40068
rect 16436 40012 20860 40068
rect 20916 40012 20926 40068
rect 22194 40012 22204 40068
rect 22260 40012 22270 40068
rect 24882 40012 24892 40068
rect 24948 40012 25340 40068
rect 25396 40012 25406 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 22204 39956 22260 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 11890 39900 11900 39956
rect 11956 39900 12572 39956
rect 12628 39900 12638 39956
rect 15698 39900 15708 39956
rect 15764 39900 17388 39956
rect 17444 39900 17454 39956
rect 18498 39900 18508 39956
rect 18564 39900 22260 39956
rect 5394 39788 5404 39844
rect 5460 39788 17276 39844
rect 17332 39788 19292 39844
rect 19348 39788 19358 39844
rect 20076 39788 21308 39844
rect 21364 39788 21868 39844
rect 21924 39788 25340 39844
rect 25396 39788 25406 39844
rect 20076 39732 20132 39788
rect 49200 39732 49800 39760
rect 9538 39676 9548 39732
rect 9604 39676 9996 39732
rect 10052 39676 10062 39732
rect 10546 39676 10556 39732
rect 10612 39676 14028 39732
rect 14084 39676 14094 39732
rect 15026 39676 15036 39732
rect 15092 39676 15428 39732
rect 15586 39676 15596 39732
rect 15652 39676 17388 39732
rect 17444 39676 17454 39732
rect 17612 39676 20132 39732
rect 20262 39676 20300 39732
rect 20356 39676 20366 39732
rect 48066 39676 48076 39732
rect 48132 39676 49800 39732
rect 15372 39620 15428 39676
rect 17612 39620 17668 39676
rect 49200 39648 49800 39676
rect 12786 39564 12796 39620
rect 12852 39564 15148 39620
rect 15204 39564 15214 39620
rect 15372 39564 17164 39620
rect 17220 39564 17668 39620
rect 20626 39564 20636 39620
rect 20692 39564 22876 39620
rect 22932 39564 23996 39620
rect 24052 39564 24062 39620
rect 25106 39564 25116 39620
rect 25172 39564 25788 39620
rect 25844 39564 25854 39620
rect 23996 39508 24052 39564
rect 12898 39452 12908 39508
rect 12964 39452 16380 39508
rect 16436 39452 17500 39508
rect 17556 39452 17566 39508
rect 17938 39452 17948 39508
rect 18004 39452 21644 39508
rect 21700 39452 21710 39508
rect 21942 39452 21980 39508
rect 22036 39452 22204 39508
rect 22260 39452 22270 39508
rect 23996 39452 25452 39508
rect 25508 39452 25518 39508
rect 7186 39340 7196 39396
rect 7252 39340 14252 39396
rect 14308 39340 14318 39396
rect 15810 39340 15820 39396
rect 15876 39340 16828 39396
rect 16884 39340 16894 39396
rect 18386 39340 18396 39396
rect 18452 39340 24332 39396
rect 24388 39340 24398 39396
rect 15586 39228 15596 39284
rect 15652 39228 16156 39284
rect 16212 39228 16222 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 9426 39116 9436 39172
rect 9492 39116 10444 39172
rect 10500 39116 10510 39172
rect 14802 39116 14812 39172
rect 14868 39116 15484 39172
rect 15540 39116 17612 39172
rect 17668 39116 17678 39172
rect 21830 39116 21868 39172
rect 21924 39116 21934 39172
rect 5954 39004 5964 39060
rect 6020 39004 11340 39060
rect 11396 39004 14028 39060
rect 14084 39004 14094 39060
rect 16034 39004 16044 39060
rect 16100 39004 16716 39060
rect 16772 39004 16782 39060
rect 19282 39004 19292 39060
rect 19348 39004 22652 39060
rect 22708 39004 22718 39060
rect 24322 39004 24332 39060
rect 24388 39004 25004 39060
rect 25060 39004 25070 39060
rect 6738 38892 6748 38948
rect 6804 38892 16156 38948
rect 16212 38892 16222 38948
rect 17826 38892 17836 38948
rect 17892 38892 29372 38948
rect 29428 38892 29438 38948
rect 14242 38780 14252 38836
rect 14308 38780 16044 38836
rect 16100 38780 16110 38836
rect 17042 38780 17052 38836
rect 17108 38780 17724 38836
rect 17780 38780 18844 38836
rect 18900 38780 18910 38836
rect 19170 38780 19180 38836
rect 19236 38780 19964 38836
rect 20020 38780 20030 38836
rect 21410 38780 21420 38836
rect 21476 38780 22988 38836
rect 23044 38780 27020 38836
rect 27076 38780 27086 38836
rect 18498 38668 18508 38724
rect 18564 38668 19068 38724
rect 19124 38668 19134 38724
rect 19618 38668 19628 38724
rect 19684 38668 19852 38724
rect 19908 38668 19918 38724
rect 20850 38668 20860 38724
rect 20916 38668 21308 38724
rect 21364 38668 21374 38724
rect 21522 38668 21532 38724
rect 21588 38668 22764 38724
rect 22820 38668 22830 38724
rect 10098 38556 10108 38612
rect 10164 38556 10892 38612
rect 10948 38556 12012 38612
rect 12068 38556 12078 38612
rect 19954 38556 19964 38612
rect 20020 38556 21588 38612
rect 19964 38500 20020 38556
rect 19142 38444 19180 38500
rect 19236 38444 19246 38500
rect 19618 38444 19628 38500
rect 19684 38444 20020 38500
rect 20374 38444 20412 38500
rect 20468 38444 20478 38500
rect 21074 38444 21084 38500
rect 21140 38444 21150 38500
rect 200 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 21084 38388 21140 38444
rect 21532 38388 21588 38556
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 200 38332 1820 38388
rect 1876 38332 1886 38388
rect 19394 38332 19404 38388
rect 19460 38332 19964 38388
rect 20020 38332 20030 38388
rect 20178 38332 20188 38388
rect 20244 38332 20860 38388
rect 20916 38332 21140 38388
rect 21522 38332 21532 38388
rect 21588 38332 27020 38388
rect 27076 38332 27086 38388
rect 200 38304 800 38332
rect 18946 38220 18956 38276
rect 19012 38220 20076 38276
rect 20132 38220 22428 38276
rect 22484 38220 22876 38276
rect 22932 38220 22942 38276
rect 10546 38108 10556 38164
rect 10612 38108 12684 38164
rect 12740 38108 12750 38164
rect 13010 38108 13020 38164
rect 13076 38108 15596 38164
rect 15652 38108 15662 38164
rect 17266 38108 17276 38164
rect 17332 38108 22764 38164
rect 22820 38108 22830 38164
rect 22950 38108 22988 38164
rect 23044 38108 23054 38164
rect 16706 37996 16716 38052
rect 16772 37996 23436 38052
rect 23492 37996 23502 38052
rect 6402 37884 6412 37940
rect 6468 37884 14812 37940
rect 14868 37884 14878 37940
rect 19170 37884 19180 37940
rect 19236 37884 20188 37940
rect 20244 37884 20254 37940
rect 20402 37884 20412 37940
rect 20468 37884 23212 37940
rect 23268 37884 23278 37940
rect 17938 37772 17948 37828
rect 18004 37772 18732 37828
rect 18788 37772 18798 37828
rect 19170 37772 19180 37828
rect 19236 37772 20300 37828
rect 20356 37772 20366 37828
rect 21746 37772 21756 37828
rect 21812 37772 22092 37828
rect 22148 37772 22158 37828
rect 49200 37716 49800 37744
rect 11554 37660 11564 37716
rect 11620 37660 19068 37716
rect 19124 37660 19134 37716
rect 19282 37660 19292 37716
rect 19348 37660 19628 37716
rect 19684 37660 19694 37716
rect 20178 37660 20188 37716
rect 20244 37660 24780 37716
rect 24836 37660 24846 37716
rect 48066 37660 48076 37716
rect 48132 37660 49800 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 49200 37632 49800 37660
rect 19142 37548 19180 37604
rect 19236 37548 19404 37604
rect 19460 37548 19470 37604
rect 11442 37436 11452 37492
rect 11508 37436 14588 37492
rect 14644 37436 15484 37492
rect 15540 37436 15550 37492
rect 18060 37436 18508 37492
rect 18564 37436 18574 37492
rect 20066 37436 20076 37492
rect 20132 37436 20972 37492
rect 21028 37436 21038 37492
rect 22502 37436 22540 37492
rect 22596 37436 22606 37492
rect 22978 37436 22988 37492
rect 23044 37436 24892 37492
rect 24948 37436 24958 37492
rect 18060 37380 18116 37436
rect 10434 37324 10444 37380
rect 10500 37324 18116 37380
rect 18274 37324 18284 37380
rect 18340 37324 20524 37380
rect 20580 37324 20590 37380
rect 20850 37324 20860 37380
rect 20916 37324 20926 37380
rect 20860 37268 20916 37324
rect 8530 37212 8540 37268
rect 8596 37212 15484 37268
rect 15540 37212 16604 37268
rect 16660 37212 20916 37268
rect 12674 37100 12684 37156
rect 12740 37100 14924 37156
rect 14980 37100 15932 37156
rect 15988 37100 15998 37156
rect 18498 37100 18508 37156
rect 18564 37100 19068 37156
rect 19124 37100 19134 37156
rect 19730 37100 19740 37156
rect 19796 37100 20300 37156
rect 20356 37100 20972 37156
rect 21028 37100 21038 37156
rect 200 37044 800 37072
rect 200 36988 1820 37044
rect 1876 36988 1886 37044
rect 16034 36988 16044 37044
rect 16100 36988 16716 37044
rect 16772 36988 16782 37044
rect 18946 36988 18956 37044
rect 19012 36988 19516 37044
rect 19572 36988 19582 37044
rect 20514 36988 20524 37044
rect 20580 36988 20860 37044
rect 20916 36988 26572 37044
rect 26628 36988 26638 37044
rect 200 36960 800 36988
rect 9090 36876 9100 36932
rect 9156 36876 15260 36932
rect 15316 36876 15326 36932
rect 15922 36876 15932 36932
rect 15988 36876 22092 36932
rect 22148 36876 22158 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 11106 36764 11116 36820
rect 11172 36764 17500 36820
rect 17556 36764 20860 36820
rect 20916 36764 23772 36820
rect 23828 36764 23838 36820
rect 26852 36764 27916 36820
rect 27972 36764 27982 36820
rect 26852 36708 26908 36764
rect 14354 36652 14364 36708
rect 14420 36652 15092 36708
rect 15148 36652 15158 36708
rect 15250 36652 15260 36708
rect 15316 36652 16156 36708
rect 16212 36652 16828 36708
rect 16884 36652 26908 36708
rect 13906 36540 13916 36596
rect 13972 36540 15036 36596
rect 15092 36540 27468 36596
rect 27524 36540 27534 36596
rect 15138 36428 15148 36484
rect 15204 36428 15242 36484
rect 15586 36428 15596 36484
rect 15652 36428 16716 36484
rect 16772 36428 18396 36484
rect 18452 36428 18462 36484
rect 19170 36428 19180 36484
rect 19236 36428 25228 36484
rect 25284 36428 25294 36484
rect 17602 36316 17612 36372
rect 17668 36316 18620 36372
rect 18676 36316 18686 36372
rect 18844 36316 24668 36372
rect 24724 36316 24734 36372
rect 18844 36260 18900 36316
rect 13682 36204 13692 36260
rect 13748 36204 14588 36260
rect 14644 36204 18900 36260
rect 19954 36204 19964 36260
rect 20020 36204 20412 36260
rect 20468 36204 20478 36260
rect 5842 36092 5852 36148
rect 5908 36092 12124 36148
rect 12180 36092 12190 36148
rect 17266 36092 17276 36148
rect 17332 36092 18060 36148
rect 18116 36092 18126 36148
rect 18274 36092 18284 36148
rect 18340 36092 19180 36148
rect 19236 36092 19246 36148
rect 18284 36036 18340 36092
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 14690 35980 14700 36036
rect 14756 35980 15148 36036
rect 15250 35980 15260 36036
rect 15316 35980 18340 36036
rect 15092 35812 15148 35980
rect 18610 35868 18620 35924
rect 18676 35868 21420 35924
rect 21476 35868 21486 35924
rect 15092 35756 26796 35812
rect 26852 35756 26862 35812
rect 49200 35700 49800 35728
rect 16594 35644 16604 35700
rect 16660 35644 21196 35700
rect 21252 35644 21262 35700
rect 48066 35644 48076 35700
rect 48132 35644 49800 35700
rect 49200 35616 49800 35644
rect 11218 35532 11228 35588
rect 11284 35532 11788 35588
rect 11844 35532 11854 35588
rect 17938 35532 17948 35588
rect 18004 35532 22540 35588
rect 22596 35532 22606 35588
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 15698 35196 15708 35252
rect 15764 35196 26236 35252
rect 26292 35196 26302 35252
rect 200 35028 800 35056
rect 200 34972 1820 35028
rect 1876 34972 1886 35028
rect 17490 34972 17500 35028
rect 17556 34972 21868 35028
rect 21924 34972 21934 35028
rect 200 34944 800 34972
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 49200 34356 49800 34384
rect 48066 34300 48076 34356
rect 48132 34300 49800 34356
rect 49200 34272 49800 34300
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 8306 33516 8316 33572
rect 8372 33516 19628 33572
rect 19684 33516 19694 33572
rect 200 33012 800 33040
rect 200 32956 1820 33012
rect 1876 32956 1886 33012
rect 200 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 49200 32340 49800 32368
rect 48066 32284 48076 32340
rect 48132 32284 49800 32340
rect 49200 32256 49800 32284
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 200 31584 800 31696
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 49200 30996 49800 31024
rect 48066 30940 48076 30996
rect 48132 30940 49800 30996
rect 49200 30912 49800 30940
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 200 29652 800 29680
rect 200 29596 1820 29652
rect 1876 29596 1886 29652
rect 200 29568 800 29596
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 49200 28980 49800 29008
rect 48066 28924 48076 28980
rect 48132 28924 49800 28980
rect 49200 28896 49800 28924
rect 200 28308 800 28336
rect 200 28252 1820 28308
rect 1876 28252 1886 28308
rect 200 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 49200 26964 49800 26992
rect 48076 26908 49800 26964
rect 48076 26852 48132 26908
rect 49200 26880 49800 26908
rect 48066 26796 48076 26852
rect 48132 26796 48142 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 200 26292 800 26320
rect 200 26236 1820 26292
rect 1876 26236 1886 26292
rect 200 26208 800 26236
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 49200 25536 49800 25648
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 200 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 200 24220 1820 24276
rect 1876 24220 1886 24276
rect 200 24192 800 24220
rect 49200 23604 49800 23632
rect 48066 23548 48076 23604
rect 48132 23548 49800 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 49200 23520 49800 23548
rect 3042 23324 3052 23380
rect 3108 23324 3500 23380
rect 3556 23324 11228 23380
rect 11284 23324 11294 23380
rect 200 22932 800 22960
rect 200 22876 2044 22932
rect 2100 22876 2110 22932
rect 200 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 49200 21588 49800 21616
rect 48066 21532 48076 21588
rect 48132 21532 49800 21588
rect 49200 21504 49800 21532
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 200 20916 800 20944
rect 200 20860 1820 20916
rect 1876 20860 1886 20916
rect 200 20832 800 20860
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 49200 20160 49800 20272
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 200 18900 800 18928
rect 200 18844 1820 18900
rect 1876 18844 1886 18900
rect 200 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 48066 18508 48076 18564
rect 48132 18508 48142 18564
rect 48076 18228 48132 18508
rect 49200 18228 49800 18256
rect 48076 18172 49800 18228
rect 49200 18144 49800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 200 17556 800 17584
rect 200 17500 1820 17556
rect 1876 17500 1886 17556
rect 200 17472 800 17500
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 49200 16884 49800 16912
rect 48066 16828 48076 16884
rect 48132 16828 49800 16884
rect 49200 16800 49800 16828
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 200 15540 800 15568
rect 200 15484 1820 15540
rect 1876 15484 1886 15540
rect 200 15456 800 15484
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 49200 14784 49800 14896
rect 200 14196 800 14224
rect 200 14140 1820 14196
rect 1876 14140 1886 14196
rect 200 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 49200 12852 49800 12880
rect 48066 12796 48076 12852
rect 48132 12796 49800 12852
rect 49200 12768 49800 12796
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 200 12096 800 12208
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 49200 11508 49800 11536
rect 48066 11452 48076 11508
rect 48132 11452 49800 11508
rect 49200 11424 49800 11452
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 200 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 200 10108 1820 10164
rect 1876 10108 1886 10164
rect 200 10080 800 10108
rect 49200 9492 49800 9520
rect 48066 9436 48076 9492
rect 48132 9436 49800 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 49200 9408 49800 9436
rect 200 8820 800 8848
rect 200 8764 1820 8820
rect 1876 8764 1886 8820
rect 200 8736 800 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 49200 7476 49800 7504
rect 48066 7420 48076 7476
rect 48132 7420 49800 7476
rect 49200 7392 49800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 200 6804 800 6832
rect 200 6748 1820 6804
rect 1876 6748 1886 6804
rect 200 6720 800 6748
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 49200 6132 49800 6160
rect 48066 6076 48076 6132
rect 48132 6076 49800 6132
rect 49200 6048 49800 6076
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 200 4704 800 4816
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 49200 4032 49800 4144
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 3042 3612 3052 3668
rect 3108 3612 4284 3668
rect 4340 3612 5852 3668
rect 5908 3612 5918 3668
rect 1362 3500 1372 3556
rect 1428 3500 2156 3556
rect 2212 3500 2222 3556
rect 200 3444 800 3472
rect 200 3388 1820 3444
rect 1876 3388 1886 3444
rect 200 3360 800 3388
rect 4722 3276 4732 3332
rect 4788 3276 5740 3332
rect 5796 3276 5806 3332
rect 28242 3276 28252 3332
rect 28308 3276 29260 3332
rect 29316 3276 29326 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 18 2268 28 2324
rect 84 2268 2492 2324
rect 2548 2268 2558 2324
rect 49200 2100 49800 2128
rect 47394 2044 47404 2100
rect 47460 2044 49800 2100
rect 49200 2016 49800 2044
rect 200 1344 800 1456
rect 49200 756 49800 784
rect 48066 700 48076 756
rect 48132 700 49800 756
rect 49200 672 49800 700
<< via3 >>
rect 14140 46284 14196 46340
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 12572 45948 12628 46004
rect 8092 45724 8148 45780
rect 10892 45724 10948 45780
rect 11004 45500 11060 45556
rect 12572 45500 12628 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 10108 45052 10164 45108
rect 16380 45052 16436 45108
rect 22540 44716 22596 44772
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 8876 44604 8932 44660
rect 21756 44604 21812 44660
rect 17052 44268 17108 44324
rect 26796 44268 26852 44324
rect 26908 44044 26964 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 21644 43708 21700 43764
rect 9100 43596 9156 43652
rect 16940 43596 16996 43652
rect 8876 43372 8932 43428
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 21868 43036 21924 43092
rect 26796 43036 26852 43092
rect 10108 42700 10164 42756
rect 26796 42700 26852 42756
rect 8316 42588 8372 42644
rect 25564 42588 25620 42644
rect 20860 42476 20916 42532
rect 25004 42476 25060 42532
rect 21980 42364 22036 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 20300 42252 20356 42308
rect 8316 42140 8372 42196
rect 14588 41804 14644 41860
rect 26684 41692 26740 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 14924 41356 14980 41412
rect 8092 41244 8148 41300
rect 10108 41132 10164 41188
rect 21756 41132 21812 41188
rect 22988 41132 23044 41188
rect 25564 41132 25620 41188
rect 19628 41020 19684 41076
rect 14140 40908 14196 40964
rect 17052 40796 17108 40852
rect 21644 40796 21700 40852
rect 22540 40796 22596 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 19404 40684 19460 40740
rect 22876 40684 22932 40740
rect 16940 40460 16996 40516
rect 14924 40348 14980 40404
rect 19180 40348 19236 40404
rect 20972 40348 21028 40404
rect 20412 40236 20468 40292
rect 26684 40236 26740 40292
rect 16380 40012 16436 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 20300 39676 20356 39732
rect 22876 39564 22932 39620
rect 21980 39452 22036 39508
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 21868 39116 21924 39172
rect 25004 39004 25060 39060
rect 19628 38668 19684 38724
rect 19180 38444 19236 38500
rect 20412 38444 20468 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19404 38332 19460 38388
rect 22988 38108 23044 38164
rect 19180 37884 19236 37940
rect 20188 37884 20244 37940
rect 20188 37660 20244 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 19180 37548 19236 37604
rect 22540 37436 22596 37492
rect 20972 37100 21028 37156
rect 9100 36876 9156 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 20860 36764 20916 36820
rect 15092 36652 15148 36708
rect 15148 36428 15204 36484
rect 14588 36204 14644 36260
rect 20412 36204 20468 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 8316 33516 8372 33572
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 14140 46340 14196 46350
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 12572 46004 12628 46014
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 8092 45780 8148 45790
rect 8092 41300 8148 45724
rect 10892 45780 10948 45790
rect 10948 45724 11060 45780
rect 10892 45714 10948 45724
rect 11004 45556 11060 45724
rect 11004 45490 11060 45500
rect 12572 45556 12628 45948
rect 12572 45490 12628 45500
rect 10108 45108 10164 45118
rect 8876 44660 8932 44670
rect 8876 43428 8932 44604
rect 8876 43362 8932 43372
rect 9100 43652 9156 43662
rect 8092 41234 8148 41244
rect 8316 42644 8372 42654
rect 8316 42196 8372 42588
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 8316 33572 8372 42140
rect 9100 36932 9156 43596
rect 10108 42756 10164 45052
rect 10108 41188 10164 42700
rect 10108 41122 10164 41132
rect 14140 40964 14196 46284
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 16380 45108 16436 45118
rect 14140 40898 14196 40908
rect 14588 41860 14644 41870
rect 9100 36866 9156 36876
rect 14588 36260 14644 41804
rect 14924 41412 14980 41422
rect 14924 40404 14980 41356
rect 14924 40338 14980 40348
rect 16380 40068 16436 45052
rect 17052 44324 17108 44334
rect 16940 43652 16996 43662
rect 16940 40516 16996 43596
rect 17052 40852 17108 44268
rect 19808 43932 20128 45444
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 22540 44772 22596 44782
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 21756 44660 21812 44670
rect 21644 43764 21700 43774
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 20860 42532 20916 42542
rect 17052 40786 17108 40796
rect 19628 41076 19684 41086
rect 16940 40450 16996 40460
rect 19404 40740 19460 40750
rect 16380 40002 16436 40012
rect 19180 40404 19236 40414
rect 19180 38500 19236 40348
rect 19180 38434 19236 38444
rect 19404 38388 19460 40684
rect 19628 38724 19684 41020
rect 19628 38658 19684 38668
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 20300 42308 20356 42318
rect 20300 39732 20356 42252
rect 20300 39666 20356 39676
rect 20412 40292 20468 40302
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19404 38322 19460 38332
rect 19180 37940 19236 37950
rect 19180 37604 19236 37884
rect 19180 37538 19236 37548
rect 19808 37660 20128 39172
rect 20412 38500 20468 40236
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 20188 37940 20244 37950
rect 20188 37716 20244 37884
rect 20188 37650 20244 37660
rect 15092 36708 15148 36718
rect 15148 36652 15204 36708
rect 15092 36642 15204 36652
rect 15148 36484 15204 36642
rect 15148 36418 15204 36428
rect 14588 36194 14644 36204
rect 8316 33506 8372 33516
rect 19808 36092 20128 37604
rect 20412 36260 20468 38444
rect 20860 36820 20916 42476
rect 21644 40852 21700 43708
rect 21756 41188 21812 44604
rect 21756 41122 21812 41132
rect 21868 43092 21924 43102
rect 21644 40786 21700 40796
rect 20972 40404 21028 40414
rect 20972 37156 21028 40348
rect 21868 39172 21924 43036
rect 21980 42420 22036 42430
rect 21980 39508 22036 42364
rect 21980 39442 22036 39452
rect 22540 40852 22596 44716
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 26796 44324 26852 44334
rect 26796 44100 26852 44268
rect 26908 44100 26964 44110
rect 26796 44044 26908 44100
rect 26908 44034 26964 44044
rect 35168 43148 35488 44660
rect 26796 43092 26852 43102
rect 26796 42756 26852 43036
rect 26796 42690 26852 42700
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 25564 42644 25620 42654
rect 25004 42532 25060 42542
rect 21868 39106 21924 39116
rect 22540 37492 22596 40796
rect 22988 41188 23044 41198
rect 22876 40740 22932 40750
rect 22876 39620 22932 40684
rect 22876 39554 22932 39564
rect 22988 38164 23044 41132
rect 25004 39060 25060 42476
rect 25564 41188 25620 42588
rect 25564 41122 25620 41132
rect 26684 41748 26740 41758
rect 26684 40292 26740 41692
rect 26684 40226 26740 40236
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 25004 38994 25060 39004
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 22988 38098 23044 38108
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 22540 37426 22596 37436
rect 20972 37090 21028 37100
rect 20860 36754 20916 36764
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 20412 36194 20468 36204
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 9072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__051__I
timestamp 1663859327
transform 1 0 23520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__052__I
timestamp 1663859327
transform -1 0 7392 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I
timestamp 1663859327
transform -1 0 7392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__054__I
timestamp 1663859327
transform 1 0 26208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__056__I
timestamp 1663859327
transform -1 0 3584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I
timestamp 1663859327
transform 1 0 20832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__058__I
timestamp 1663859327
transform 1 0 13104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I
timestamp 1663859327
transform 1 0 14896 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__060__I
timestamp 1663859327
transform 1 0 29792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__061__I
timestamp 1663859327
transform 1 0 22400 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I
timestamp 1663859327
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I
timestamp 1663859327
transform 1 0 20272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__065__I
timestamp 1663859327
transform 1 0 27552 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I
timestamp 1663859327
transform 1 0 30352 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__067__I
timestamp 1663859327
transform -1 0 17136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I
timestamp 1663859327
transform -1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__069__I
timestamp 1663859327
transform -1 0 5376 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__070__I
timestamp 1663859327
transform -1 0 7840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I
timestamp 1663859327
transform -1 0 25424 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__072__I
timestamp 1663859327
transform 1 0 18928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I
timestamp 1663859327
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__074__I
timestamp 1663859327
transform -1 0 22176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I
timestamp 1663859327
transform 1 0 4480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__A1
timestamp 1663859327
transform -1 0 16240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__076__A2
timestamp 1663859327
transform 1 0 14224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I
timestamp 1663859327
transform 1 0 26656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__A1
timestamp 1663859327
transform -1 0 5152 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__078__A2
timestamp 1663859327
transform -1 0 4032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__A1
timestamp 1663859327
transform 1 0 26656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__A2
timestamp 1663859327
transform 1 0 25760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__A3
timestamp 1663859327
transform 1 0 26208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__A1
timestamp 1663859327
transform -1 0 18704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__B
timestamp 1663859327
transform -1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I
timestamp 1663859327
transform 1 0 28896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__A1
timestamp 1663859327
transform 1 0 21504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__A2
timestamp 1663859327
transform 1 0 20832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__082__A3
timestamp 1663859327
transform -1 0 20048 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I
timestamp 1663859327
transform -1 0 15568 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1663859327
transform -1 0 6272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__A1
timestamp 1663859327
transform 1 0 7392 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__A2
timestamp 1663859327
transform -1 0 4704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__A3
timestamp 1663859327
transform 1 0 8064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__A4
timestamp 1663859327
transform 1 0 5152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__086__A1
timestamp 1663859327
transform 1 0 10192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__A1
timestamp 1663859327
transform 1 0 27552 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__A2
timestamp 1663859327
transform 1 0 29456 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__B
timestamp 1663859327
transform 1 0 30352 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__A1
timestamp 1663859327
transform -1 0 18256 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__088__A2
timestamp 1663859327
transform -1 0 18704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__A1
timestamp 1663859327
transform 1 0 10976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__A2
timestamp 1663859327
transform 1 0 10528 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__B
timestamp 1663859327
transform 1 0 9968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I
timestamp 1663859327
transform 1 0 19376 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__A1
timestamp 1663859327
transform -1 0 9968 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__A2
timestamp 1663859327
transform -1 0 11088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__091__C
timestamp 1663859327
transform 1 0 8288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__A1
timestamp 1663859327
transform -1 0 19152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__A2
timestamp 1663859327
transform -1 0 20944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__A1
timestamp 1663859327
transform -1 0 5040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__A2
timestamp 1663859327
transform -1 0 19152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__A3
timestamp 1663859327
transform -1 0 4592 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__093__A4
timestamp 1663859327
transform -1 0 4144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__A1
timestamp 1663859327
transform -1 0 20944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A1
timestamp 1663859327
transform 1 0 24416 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A2
timestamp 1663859327
transform 1 0 23968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__095__A3
timestamp 1663859327
transform -1 0 23072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__A1
timestamp 1663859327
transform 1 0 27104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__097__B
timestamp 1663859327
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__A1
timestamp 1663859327
transform 1 0 15120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__A2
timestamp 1663859327
transform -1 0 14224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I
timestamp 1663859327
transform -1 0 11984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__100__I
timestamp 1663859327
transform 1 0 30800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A1
timestamp 1663859327
transform -1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A2
timestamp 1663859327
transform -1 0 17808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__A3
timestamp 1663859327
transform -1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A1
timestamp 1663859327
transform 1 0 29344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__A2
timestamp 1663859327
transform 1 0 28000 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__A1
timestamp 1663859327
transform 1 0 10640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__A2
timestamp 1663859327
transform -1 0 11536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__B
timestamp 1663859327
transform -1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A1
timestamp 1663859327
transform 1 0 5600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__104__A2
timestamp 1663859327
transform -1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A1
timestamp 1663859327
transform -1 0 8288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__A2
timestamp 1663859327
transform 1 0 10416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__A1
timestamp 1663859327
transform -1 0 4928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__A2
timestamp 1663859327
transform -1 0 3808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__106__B2
timestamp 1663859327
transform -1 0 8848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A1
timestamp 1663859327
transform 1 0 32144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__A2
timestamp 1663859327
transform 1 0 29904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__B
timestamp 1663859327
transform 1 0 29344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A1
timestamp 1663859327
transform 1 0 25312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A2
timestamp 1663859327
transform 1 0 22064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__A2
timestamp 1663859327
transform 1 0 23744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__109__C
timestamp 1663859327
transform 1 0 26880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__A1
timestamp 1663859327
transform 1 0 28448 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__A1
timestamp 1663859327
transform -1 0 23072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__A2
timestamp 1663859327
transform 1 0 23744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__A1
timestamp 1663859327
transform 1 0 28000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A1
timestamp 1663859327
transform 1 0 31136 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A2
timestamp 1663859327
transform 1 0 31248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__B
timestamp 1663859327
transform 1 0 31584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__A1
timestamp 1663859327
transform -1 0 9184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__A2
timestamp 1663859327
transform -1 0 13776 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__B1
timestamp 1663859327
transform -1 0 10640 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__B2
timestamp 1663859327
transform 1 0 7840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__A1
timestamp 1663859327
transform -1 0 25088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__A2
timestamp 1663859327
transform -1 0 27328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__A1
timestamp 1663859327
transform -1 0 12432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__A2
timestamp 1663859327
transform 1 0 15568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__B
timestamp 1663859327
transform -1 0 12880 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__A1
timestamp 1663859327
transform -1 0 24416 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__A2
timestamp 1663859327
transform -1 0 27776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__B2
timestamp 1663859327
transform 1 0 26208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__A1
timestamp 1663859327
transform -1 0 8736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__A2
timestamp 1663859327
transform -1 0 14784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__A3
timestamp 1663859327
transform -1 0 7840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__A1
timestamp 1663859327
transform 1 0 23072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__A2
timestamp 1663859327
transform 1 0 23296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__A3
timestamp 1663859327
transform 1 0 22400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__A1
timestamp 1663859327
transform -1 0 20496 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__A2
timestamp 1663859327
transform -1 0 19600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__A1
timestamp 1663859327
transform -1 0 21840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__A2
timestamp 1663859327
transform 1 0 21168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__B
timestamp 1663859327
transform -1 0 20496 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__A1
timestamp 1663859327
transform 1 0 30688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__A2
timestamp 1663859327
transform 1 0 32032 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__B
timestamp 1663859327
transform 1 0 29456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1663859327
transform -1 0 14000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A1
timestamp 1663859327
transform 1 0 28896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A2
timestamp 1663859327
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__A1
timestamp 1663859327
transform 1 0 9632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__A2
timestamp 1663859327
transform -1 0 9632 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1663859327
transform 1 0 31136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A1
timestamp 1663859327
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A2
timestamp 1663859327
transform 1 0 31696 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__B
timestamp 1663859327
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__CLKN
timestamp 1663859327
transform 1 0 32592 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__CLKN
timestamp 1663859327
transform -1 0 18032 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__CLKN
timestamp 1663859327
transform 1 0 3472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__CLK
timestamp 1663859327
transform 1 0 28000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__D
timestamp 1663859327
transform -1 0 7168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__CLK
timestamp 1663859327
transform -1 0 7616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__D
timestamp 1663859327
transform -1 0 6272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__CLK
timestamp 1663859327
transform 1 0 22960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__D
timestamp 1663859327
transform 1 0 25984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__CLK
timestamp 1663859327
transform 1 0 21504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__D
timestamp 1663859327
transform -1 0 20048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__CLK
timestamp 1663859327
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__D
timestamp 1663859327
transform -1 0 23520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__CLK
timestamp 1663859327
transform -1 0 22176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__D
timestamp 1663859327
transform 1 0 30240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__CLK
timestamp 1663859327
transform -1 0 16240 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__D
timestamp 1663859327
transform -1 0 17584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__CLK
timestamp 1663859327
transform -1 0 21056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__CLK
timestamp 1663859327
transform 1 0 31920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__D
timestamp 1663859327
transform 1 0 32368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__CLK
timestamp 1663859327
transform -1 0 3248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__143__D
timestamp 1663859327
transform -1 0 4256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__CLK
timestamp 1663859327
transform -1 0 6720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__D
timestamp 1663859327
transform -1 0 5824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__CLK
timestamp 1663859327
transform -1 0 14672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__CLK
timestamp 1663859327
transform 1 0 6720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__CLK
timestamp 1663859327
transform -1 0 12656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__D
timestamp 1663859327
transform 1 0 11312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__148__CLK
timestamp 1663859327
transform 1 0 11984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__CLK
timestamp 1663859327
transform 1 0 25760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__CLK
timestamp 1663859327
transform -1 0 6272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__D
timestamp 1663859327
transform -1 0 6720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__CLKN
timestamp 1663859327
transform 1 0 27328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__CLK
timestamp 1663859327
transform 1 0 9968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__D
timestamp 1663859327
transform -1 0 7168 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__CLK
timestamp 1663859327
transform -1 0 1904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__D
timestamp 1663859327
transform -1 0 6496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__CLK
timestamp 1663859327
transform 1 0 5600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__D
timestamp 1663859327
transform -1 0 8400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__CLK
timestamp 1663859327
transform 1 0 22512 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__CLKN
timestamp 1663859327
transform 1 0 9520 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__CLKN
timestamp 1663859327
transform 1 0 10864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__CLKN
timestamp 1663859327
transform 1 0 4256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1663859327
transform -1 0 8736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1663859327
transform 1 0 31584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output5_I
timestamp 1663859327
transform 1 0 34720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output6_I
timestamp 1663859327
transform -1 0 3136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output7_I
timestamp 1663859327
transform 1 0 3472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1663859327
transform -1 0 4368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output9_I
timestamp 1663859327
transform -1 0 42560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1663859327
transform 1 0 33488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 3248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23
timestamp 1663859327
transform 1 0 3920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 4368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1663859327
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 6048 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58
timestamp 1663859327
transform 1 0 7840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1663859327
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77
timestamp 1663859327
transform 1 0 9968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93
timestamp 1663859327
transform 1 0 11760 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_101
timestamp 1663859327
transform 1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1663859327
transform 1 0 13328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119
timestamp 1663859327
transform 1 0 14672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_131
timestamp 1663859327
transform 1 0 16016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1663859327
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1663859327
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1663859327
transform 1 0 17472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_149
timestamp 1663859327
transform 1 0 18032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_165
timestamp 1663859327
transform 1 0 19824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1663859327
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1663859327
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_182
timestamp 1663859327
transform 1 0 21728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190
timestamp 1663859327
transform 1 0 22624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192
timestamp 1663859327
transform 1 0 22848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_197
timestamp 1663859327
transform 1 0 23408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_205
timestamp 1663859327
transform 1 0 24304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1663859327
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_212
timestamp 1663859327
transform 1 0 25088 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1663859327
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_222
timestamp 1663859327
transform 1 0 26208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_227
timestamp 1663859327
transform 1 0 26768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_243
timestamp 1663859327
transform 1 0 28560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1663859327
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_252
timestamp 1663859327
transform 1 0 29568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_268
timestamp 1663859327
transform 1 0 31360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_270
timestamp 1663859327
transform 1 0 31584 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_275
timestamp 1663859327
transform 1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1663859327
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_282
timestamp 1663859327
transform 1 0 32928 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_298
timestamp 1663859327
transform 1 0 34720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_300
timestamp 1663859327
transform 1 0 34944 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_305
timestamp 1663859327
transform 1 0 35504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1663859327
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_317
timestamp 1663859327
transform 1 0 36848 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_325
timestamp 1663859327
transform 1 0 37744 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329
timestamp 1663859327
transform 1 0 38192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_335
timestamp 1663859327
transform 1 0 38864 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_343
timestamp 1663859327
transform 1 0 39760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1663859327
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1663859327
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1663859327
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_357
timestamp 1663859327
transform 1 0 41328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_365
timestamp 1663859327
transform 1 0 42224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_371
timestamp 1663859327
transform 1 0 42896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_383
timestamp 1663859327
transform 1 0 44240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_387
timestamp 1663859327
transform 1 0 44688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_395
timestamp 1663859327
transform 1 0 45584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_401
timestamp 1663859327
transform 1 0 46256 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_413
timestamp 1663859327
transform 1 0 47600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1663859327
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1663859327
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_7
timestamp 1663859327
transform 1 0 2128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_13 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2800 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_45
timestamp 1663859327
transform 1 0 6384 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_61
timestamp 1663859327
transform 1 0 8176 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_69
timestamp 1663859327
transform 1 0 9072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1663859327
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1663859327
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1663859327
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1663859327
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1663859327
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1663859327
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1663859327
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1663859327
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1663859327
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1663859327
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1663859327
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_357
timestamp 1663859327
transform 1 0 41328 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_389
timestamp 1663859327
transform 1 0 44912 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_405
timestamp 1663859327
transform 1 0 46704 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_413
timestamp 1663859327
transform 1 0 47600 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_417
timestamp 1663859327
transform 1 0 48048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1663859327
transform 1 0 48272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1663859327
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1663859327
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1663859327
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1663859327
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1663859327
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1663859327
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1663859327
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1663859327
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1663859327
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1663859327
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1663859327
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1663859327
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1663859327
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1663859327
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1663859327
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1663859327
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1663859327
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1663859327
transform 1 0 45248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_408
timestamp 1663859327
transform 1 0 47040 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_416
timestamp 1663859327
transform 1 0 47936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1663859327
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1663859327
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1663859327
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1663859327
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1663859327
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1663859327
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1663859327
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1663859327
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1663859327
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1663859327
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1663859327
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1663859327
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1663859327
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1663859327
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1663859327
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_357
timestamp 1663859327
transform 1 0 41328 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_389
timestamp 1663859327
transform 1 0 44912 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_405
timestamp 1663859327
transform 1 0 46704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1663859327
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1663859327
transform 1 0 48048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1663859327
transform 1 0 48272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1663859327
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1663859327
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1663859327
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1663859327
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1663859327
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1663859327
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1663859327
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1663859327
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1663859327
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1663859327
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1663859327
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1663859327
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1663859327
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1663859327
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1663859327
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1663859327
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1663859327
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_392
timestamp 1663859327
transform 1 0 45248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_408
timestamp 1663859327
transform 1 0 47040 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_412
timestamp 1663859327
transform 1 0 47488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_414
timestamp 1663859327
transform 1 0 47712 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_419
timestamp 1663859327
transform 1 0 48272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1663859327
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_7
timestamp 1663859327
transform 1 0 2128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1663859327
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1663859327
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1663859327
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1663859327
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1663859327
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1663859327
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1663859327
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1663859327
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1663859327
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1663859327
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1663859327
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1663859327
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_357
timestamp 1663859327
transform 1 0 41328 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_389
timestamp 1663859327
transform 1 0 44912 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_405
timestamp 1663859327
transform 1 0 46704 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1663859327
transform 1 0 47600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1663859327
transform 1 0 48048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1663859327
transform 1 0 48272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1663859327
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1663859327
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1663859327
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1663859327
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1663859327
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1663859327
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1663859327
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1663859327
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1663859327
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1663859327
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1663859327
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1663859327
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1663859327
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1663859327
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1663859327
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1663859327
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1663859327
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_392
timestamp 1663859327
transform 1 0 45248 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_408
timestamp 1663859327
transform 1 0 47040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_412
timestamp 1663859327
transform 1 0 47488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_414
timestamp 1663859327
transform 1 0 47712 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1663859327
transform 1 0 48272 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1663859327
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_7
timestamp 1663859327
transform 1 0 2128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1663859327
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1663859327
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1663859327
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1663859327
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1663859327
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1663859327
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1663859327
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1663859327
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1663859327
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1663859327
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1663859327
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1663859327
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_357
timestamp 1663859327
transform 1 0 41328 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_389
timestamp 1663859327
transform 1 0 44912 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_405
timestamp 1663859327
transform 1 0 46704 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_413
timestamp 1663859327
transform 1 0 47600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1663859327
transform 1 0 48048 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1663859327
transform 1 0 48272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1663859327
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1663859327
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1663859327
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1663859327
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1663859327
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1663859327
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1663859327
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1663859327
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1663859327
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1663859327
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1663859327
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1663859327
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1663859327
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1663859327
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1663859327
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1663859327
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1663859327
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_392
timestamp 1663859327
transform 1 0 45248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_408
timestamp 1663859327
transform 1 0 47040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_412
timestamp 1663859327
transform 1 0 47488 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_414
timestamp 1663859327
transform 1 0 47712 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_419
timestamp 1663859327
transform 1 0 48272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1663859327
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_7
timestamp 1663859327
transform 1 0 2128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1663859327
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1663859327
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1663859327
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1663859327
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1663859327
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1663859327
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1663859327
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1663859327
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1663859327
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1663859327
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1663859327
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1663859327
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_357
timestamp 1663859327
transform 1 0 41328 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_389
timestamp 1663859327
transform 1 0 44912 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1663859327
transform 1 0 46704 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1663859327
transform 1 0 47600 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1663859327
transform 1 0 48048 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1663859327
transform 1 0 48272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1663859327
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1663859327
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1663859327
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1663859327
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1663859327
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1663859327
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1663859327
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1663859327
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1663859327
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1663859327
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1663859327
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1663859327
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1663859327
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1663859327
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1663859327
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1663859327
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1663859327
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1663859327
transform 1 0 45248 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1663859327
transform 1 0 47040 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1663859327
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1663859327
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1663859327
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1663859327
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1663859327
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1663859327
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1663859327
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1663859327
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1663859327
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1663859327
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1663859327
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1663859327
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1663859327
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1663859327
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1663859327
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1663859327
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_357
timestamp 1663859327
transform 1 0 41328 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_389
timestamp 1663859327
transform 1 0 44912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_405
timestamp 1663859327
transform 1 0 46704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_413
timestamp 1663859327
transform 1 0 47600 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1663859327
transform 1 0 48272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1663859327
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1663859327
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1663859327
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1663859327
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1663859327
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1663859327
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1663859327
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1663859327
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1663859327
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1663859327
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1663859327
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1663859327
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1663859327
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1663859327
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1663859327
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1663859327
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1663859327
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_392
timestamp 1663859327
transform 1 0 45248 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_408
timestamp 1663859327
transform 1 0 47040 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_412
timestamp 1663859327
transform 1 0 47488 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_414
timestamp 1663859327
transform 1 0 47712 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_419
timestamp 1663859327
transform 1 0 48272 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1663859327
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1663859327
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1663859327
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1663859327
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1663859327
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1663859327
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1663859327
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1663859327
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1663859327
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1663859327
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1663859327
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1663859327
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1663859327
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1663859327
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1663859327
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_357
timestamp 1663859327
transform 1 0 41328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_389
timestamp 1663859327
transform 1 0 44912 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_405
timestamp 1663859327
transform 1 0 46704 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_413
timestamp 1663859327
transform 1 0 47600 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1663859327
transform 1 0 48048 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1663859327
transform 1 0 48272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1663859327
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_7
timestamp 1663859327
transform 1 0 2128 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_23
timestamp 1663859327
transform 1 0 3920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_31
timestamp 1663859327
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1663859327
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1663859327
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1663859327
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1663859327
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1663859327
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1663859327
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1663859327
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1663859327
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1663859327
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1663859327
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1663859327
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1663859327
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1663859327
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1663859327
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1663859327
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_392
timestamp 1663859327
transform 1 0 45248 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1663859327
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_416
timestamp 1663859327
transform 1 0 47936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1663859327
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1663859327
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1663859327
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1663859327
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1663859327
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1663859327
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1663859327
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1663859327
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1663859327
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1663859327
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1663859327
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1663859327
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1663859327
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1663859327
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1663859327
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_357
timestamp 1663859327
transform 1 0 41328 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_389
timestamp 1663859327
transform 1 0 44912 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_405
timestamp 1663859327
transform 1 0 46704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_413
timestamp 1663859327
transform 1 0 47600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_417
timestamp 1663859327
transform 1 0 48048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1663859327
transform 1 0 48272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1663859327
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_7
timestamp 1663859327
transform 1 0 2128 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_23
timestamp 1663859327
transform 1 0 3920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_31
timestamp 1663859327
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1663859327
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1663859327
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1663859327
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1663859327
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1663859327
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1663859327
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1663859327
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1663859327
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1663859327
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1663859327
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1663859327
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1663859327
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1663859327
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1663859327
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1663859327
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_392
timestamp 1663859327
transform 1 0 45248 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_408
timestamp 1663859327
transform 1 0 47040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_416
timestamp 1663859327
transform 1 0 47936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1663859327
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1663859327
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1663859327
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1663859327
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1663859327
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1663859327
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1663859327
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1663859327
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1663859327
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1663859327
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1663859327
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1663859327
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1663859327
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1663859327
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1663859327
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_357
timestamp 1663859327
transform 1 0 41328 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_389
timestamp 1663859327
transform 1 0 44912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_405
timestamp 1663859327
transform 1 0 46704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_413
timestamp 1663859327
transform 1 0 47600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_417
timestamp 1663859327
transform 1 0 48048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1663859327
transform 1 0 48272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1663859327
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_7
timestamp 1663859327
transform 1 0 2128 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_23
timestamp 1663859327
transform 1 0 3920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_31
timestamp 1663859327
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1663859327
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1663859327
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1663859327
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1663859327
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1663859327
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1663859327
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1663859327
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1663859327
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1663859327
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1663859327
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1663859327
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1663859327
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1663859327
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1663859327
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1663859327
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_392
timestamp 1663859327
transform 1 0 45248 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_408
timestamp 1663859327
transform 1 0 47040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_412
timestamp 1663859327
transform 1 0 47488 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_414
timestamp 1663859327
transform 1 0 47712 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_419
timestamp 1663859327
transform 1 0 48272 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1663859327
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1663859327
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1663859327
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1663859327
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1663859327
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1663859327
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1663859327
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1663859327
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1663859327
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1663859327
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1663859327
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1663859327
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1663859327
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1663859327
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1663859327
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_357
timestamp 1663859327
transform 1 0 41328 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_389
timestamp 1663859327
transform 1 0 44912 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_405
timestamp 1663859327
transform 1 0 46704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_413
timestamp 1663859327
transform 1 0 47600 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_419
timestamp 1663859327
transform 1 0 48272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_2
timestamp 1663859327
transform 1 0 1568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_7
timestamp 1663859327
transform 1 0 2128 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_23
timestamp 1663859327
transform 1 0 3920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_31
timestamp 1663859327
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1663859327
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1663859327
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1663859327
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1663859327
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1663859327
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1663859327
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1663859327
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1663859327
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1663859327
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1663859327
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1663859327
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1663859327
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1663859327
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1663859327
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1663859327
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_392
timestamp 1663859327
transform 1 0 45248 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_408
timestamp 1663859327
transform 1 0 47040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_416
timestamp 1663859327
transform 1 0 47936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1663859327
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1663859327
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1663859327
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1663859327
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1663859327
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1663859327
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1663859327
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1663859327
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1663859327
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1663859327
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1663859327
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1663859327
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1663859327
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1663859327
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1663859327
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_357
timestamp 1663859327
transform 1 0 41328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_389
timestamp 1663859327
transform 1 0 44912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_405
timestamp 1663859327
transform 1 0 46704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_413
timestamp 1663859327
transform 1 0 47600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_417
timestamp 1663859327
transform 1 0 48048 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_419
timestamp 1663859327
transform 1 0 48272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1663859327
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1663859327
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1663859327
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1663859327
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1663859327
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1663859327
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1663859327
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1663859327
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1663859327
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1663859327
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1663859327
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1663859327
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1663859327
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1663859327
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1663859327
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1663859327
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1663859327
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_392
timestamp 1663859327
transform 1 0 45248 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_408
timestamp 1663859327
transform 1 0 47040 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_416
timestamp 1663859327
transform 1 0 47936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1663859327
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_7
timestamp 1663859327
transform 1 0 2128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1663859327
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1663859327
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1663859327
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1663859327
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1663859327
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1663859327
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1663859327
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1663859327
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1663859327
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1663859327
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1663859327
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1663859327
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_357
timestamp 1663859327
transform 1 0 41328 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_389
timestamp 1663859327
transform 1 0 44912 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_405
timestamp 1663859327
transform 1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_413
timestamp 1663859327
transform 1 0 47600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_417
timestamp 1663859327
transform 1 0 48048 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_419
timestamp 1663859327
transform 1 0 48272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1663859327
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1663859327
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1663859327
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1663859327
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1663859327
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1663859327
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1663859327
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1663859327
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1663859327
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1663859327
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1663859327
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1663859327
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1663859327
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1663859327
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1663859327
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1663859327
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1663859327
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_392
timestamp 1663859327
transform 1 0 45248 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_408
timestamp 1663859327
transform 1 0 47040 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_412
timestamp 1663859327
transform 1 0 47488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_414
timestamp 1663859327
transform 1 0 47712 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_419
timestamp 1663859327
transform 1 0 48272 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1663859327
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_17
timestamp 1663859327
transform 1 0 3248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_21
timestamp 1663859327
transform 1 0 3696 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_53
timestamp 1663859327
transform 1 0 7280 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_69
timestamp 1663859327
transform 1 0 9072 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1663859327
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1663859327
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1663859327
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1663859327
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1663859327
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1663859327
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1663859327
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1663859327
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1663859327
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1663859327
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1663859327
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1663859327
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_357
timestamp 1663859327
transform 1 0 41328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_389
timestamp 1663859327
transform 1 0 44912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_405
timestamp 1663859327
transform 1 0 46704 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_413
timestamp 1663859327
transform 1 0 47600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_417
timestamp 1663859327
transform 1 0 48048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_419
timestamp 1663859327
transform 1 0 48272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1663859327
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1663859327
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1663859327
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1663859327
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1663859327
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1663859327
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1663859327
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1663859327
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1663859327
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1663859327
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1663859327
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1663859327
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1663859327
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1663859327
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1663859327
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1663859327
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1663859327
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_392
timestamp 1663859327
transform 1 0 45248 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_408
timestamp 1663859327
transform 1 0 47040 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_412
timestamp 1663859327
transform 1 0 47488 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_414
timestamp 1663859327
transform 1 0 47712 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_419
timestamp 1663859327
transform 1 0 48272 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1663859327
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_7
timestamp 1663859327
transform 1 0 2128 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1663859327
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1663859327
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1663859327
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1663859327
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1663859327
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1663859327
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1663859327
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1663859327
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1663859327
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1663859327
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1663859327
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1663859327
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_357
timestamp 1663859327
transform 1 0 41328 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_389
timestamp 1663859327
transform 1 0 44912 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_405
timestamp 1663859327
transform 1 0 46704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_413
timestamp 1663859327
transform 1 0 47600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_417
timestamp 1663859327
transform 1 0 48048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1663859327
transform 1 0 48272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1663859327
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1663859327
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1663859327
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1663859327
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1663859327
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1663859327
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1663859327
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1663859327
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1663859327
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1663859327
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1663859327
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1663859327
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1663859327
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1663859327
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1663859327
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1663859327
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1663859327
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_392
timestamp 1663859327
transform 1 0 45248 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_408
timestamp 1663859327
transform 1 0 47040 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_416
timestamp 1663859327
transform 1 0 47936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1663859327
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1663859327
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1663859327
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1663859327
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1663859327
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1663859327
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1663859327
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1663859327
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1663859327
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1663859327
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1663859327
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1663859327
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1663859327
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1663859327
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1663859327
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_357
timestamp 1663859327
transform 1 0 41328 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_389
timestamp 1663859327
transform 1 0 44912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_405
timestamp 1663859327
transform 1 0 46704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_413
timestamp 1663859327
transform 1 0 47600 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_417
timestamp 1663859327
transform 1 0 48048 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1663859327
transform 1 0 48272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1663859327
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_7
timestamp 1663859327
transform 1 0 2128 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_23
timestamp 1663859327
transform 1 0 3920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_31
timestamp 1663859327
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1663859327
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1663859327
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1663859327
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1663859327
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1663859327
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1663859327
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1663859327
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1663859327
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1663859327
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1663859327
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1663859327
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1663859327
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1663859327
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1663859327
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1663859327
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_392
timestamp 1663859327
transform 1 0 45248 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_408
timestamp 1663859327
transform 1 0 47040 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_412
timestamp 1663859327
transform 1 0 47488 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_414
timestamp 1663859327
transform 1 0 47712 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_419
timestamp 1663859327
transform 1 0 48272 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1663859327
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1663859327
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1663859327
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1663859327
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1663859327
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1663859327
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1663859327
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1663859327
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1663859327
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1663859327
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1663859327
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1663859327
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1663859327
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1663859327
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1663859327
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_357
timestamp 1663859327
transform 1 0 41328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_389
timestamp 1663859327
transform 1 0 44912 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_405
timestamp 1663859327
transform 1 0 46704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_413
timestamp 1663859327
transform 1 0 47600 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_417
timestamp 1663859327
transform 1 0 48048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_419
timestamp 1663859327
transform 1 0 48272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1663859327
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_7
timestamp 1663859327
transform 1 0 2128 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_23
timestamp 1663859327
transform 1 0 3920 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_31
timestamp 1663859327
transform 1 0 4816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1663859327
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1663859327
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1663859327
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1663859327
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1663859327
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1663859327
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1663859327
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1663859327
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1663859327
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1663859327
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1663859327
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1663859327
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1663859327
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1663859327
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1663859327
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_392
timestamp 1663859327
transform 1 0 45248 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_408
timestamp 1663859327
transform 1 0 47040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_416
timestamp 1663859327
transform 1 0 47936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1663859327
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1663859327
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1663859327
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1663859327
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1663859327
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1663859327
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1663859327
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1663859327
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1663859327
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1663859327
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1663859327
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1663859327
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1663859327
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1663859327
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1663859327
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_357
timestamp 1663859327
transform 1 0 41328 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_389
timestamp 1663859327
transform 1 0 44912 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_405
timestamp 1663859327
transform 1 0 46704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_413
timestamp 1663859327
transform 1 0 47600 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_419
timestamp 1663859327
transform 1 0 48272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1663859327
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_7
timestamp 1663859327
transform 1 0 2128 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_23
timestamp 1663859327
transform 1 0 3920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_31
timestamp 1663859327
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1663859327
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1663859327
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1663859327
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1663859327
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1663859327
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1663859327
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1663859327
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1663859327
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1663859327
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1663859327
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1663859327
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1663859327
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1663859327
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1663859327
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1663859327
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_392
timestamp 1663859327
transform 1 0 45248 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_408
timestamp 1663859327
transform 1 0 47040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_416
timestamp 1663859327
transform 1 0 47936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1663859327
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1663859327
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1663859327
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1663859327
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1663859327
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1663859327
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1663859327
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1663859327
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1663859327
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1663859327
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1663859327
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1663859327
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1663859327
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1663859327
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1663859327
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_357
timestamp 1663859327
transform 1 0 41328 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_389
timestamp 1663859327
transform 1 0 44912 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_405
timestamp 1663859327
transform 1 0 46704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_413
timestamp 1663859327
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_417
timestamp 1663859327
transform 1 0 48048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_419
timestamp 1663859327
transform 1 0 48272 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1663859327
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1663859327
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1663859327
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1663859327
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1663859327
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1663859327
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1663859327
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1663859327
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1663859327
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1663859327
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1663859327
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1663859327
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1663859327
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1663859327
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1663859327
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1663859327
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1663859327
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_392
timestamp 1663859327
transform 1 0 45248 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_408
timestamp 1663859327
transform 1 0 47040 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_412
timestamp 1663859327
transform 1 0 47488 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_414
timestamp 1663859327
transform 1 0 47712 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_419
timestamp 1663859327
transform 1 0 48272 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1663859327
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1663859327
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1663859327
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1663859327
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1663859327
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1663859327
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1663859327
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1663859327
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1663859327
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1663859327
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1663859327
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1663859327
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1663859327
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1663859327
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1663859327
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_357
timestamp 1663859327
transform 1 0 41328 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_389
timestamp 1663859327
transform 1 0 44912 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_405
timestamp 1663859327
transform 1 0 46704 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_413
timestamp 1663859327
transform 1 0 47600 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_419
timestamp 1663859327
transform 1 0 48272 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1663859327
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_7
timestamp 1663859327
transform 1 0 2128 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_23
timestamp 1663859327
transform 1 0 3920 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_31
timestamp 1663859327
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1663859327
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1663859327
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1663859327
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1663859327
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1663859327
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1663859327
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1663859327
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1663859327
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1663859327
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1663859327
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1663859327
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1663859327
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1663859327
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1663859327
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1663859327
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_392
timestamp 1663859327
transform 1 0 45248 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_408
timestamp 1663859327
transform 1 0 47040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_416
timestamp 1663859327
transform 1 0 47936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1663859327
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1663859327
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1663859327
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1663859327
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1663859327
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1663859327
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1663859327
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1663859327
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1663859327
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1663859327
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1663859327
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1663859327
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1663859327
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1663859327
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1663859327
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1663859327
transform 1 0 41328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_389
timestamp 1663859327
transform 1 0 44912 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_405
timestamp 1663859327
transform 1 0 46704 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_413
timestamp 1663859327
transform 1 0 47600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_417
timestamp 1663859327
transform 1 0 48048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_419
timestamp 1663859327
transform 1 0 48272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1663859327
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1663859327
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1663859327
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1663859327
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1663859327
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_108
timestamp 1663859327
transform 1 0 13440 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_140
timestamp 1663859327
transform 1 0 17024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_142
timestamp 1663859327
transform 1 0 17248 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_145
timestamp 1663859327
transform 1 0 17584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_149
timestamp 1663859327
transform 1 0 18032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_155
timestamp 1663859327
transform 1 0 18704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_159
timestamp 1663859327
transform 1 0 19152 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_175
timestamp 1663859327
transform 1 0 20944 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1663859327
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1663859327
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1663859327
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1663859327
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1663859327
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1663859327
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1663859327
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1663859327
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1663859327
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_392
timestamp 1663859327
transform 1 0 45248 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_408
timestamp 1663859327
transform 1 0 47040 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_412
timestamp 1663859327
transform 1 0 47488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_414
timestamp 1663859327
transform 1 0 47712 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_419
timestamp 1663859327
transform 1 0 48272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1663859327
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_7
timestamp 1663859327
transform 1 0 2128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_73
timestamp 1663859327
transform 1 0 9520 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_105
timestamp 1663859327
transform 1 0 13104 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_121
timestamp 1663859327
transform 1 0 14896 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_129
timestamp 1663859327
transform 1 0 15792 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_133
timestamp 1663859327
transform 1 0 16240 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_137
timestamp 1663859327
transform 1 0 16688 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1663859327
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1663859327
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_147
timestamp 1663859327
transform 1 0 17808 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_151
timestamp 1663859327
transform 1 0 18256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_155
timestamp 1663859327
transform 1 0 18704 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_159
timestamp 1663859327
transform 1 0 19152 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_163
timestamp 1663859327
transform 1 0 19600 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_167
timestamp 1663859327
transform 1 0 20048 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_171
timestamp 1663859327
transform 1 0 20496 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_175
timestamp 1663859327
transform 1 0 20944 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_207
timestamp 1663859327
transform 1 0 24528 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_211
timestamp 1663859327
transform 1 0 24976 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1663859327
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1663859327
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1663859327
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1663859327
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1663859327
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1663859327
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_357
timestamp 1663859327
transform 1 0 41328 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_389
timestamp 1663859327
transform 1 0 44912 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_405
timestamp 1663859327
transform 1 0 46704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_413
timestamp 1663859327
transform 1 0 47600 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_417
timestamp 1663859327
transform 1 0 48048 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_419
timestamp 1663859327
transform 1 0 48272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1663859327
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1663859327
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1663859327
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1663859327
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1663859327
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_108
timestamp 1663859327
transform 1 0 13440 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_116
timestamp 1663859327
transform 1 0 14336 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_120
timestamp 1663859327
transform 1 0 14784 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_122
timestamp 1663859327
transform 1 0 15008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_125
timestamp 1663859327
transform 1 0 15344 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_129
timestamp 1663859327
transform 1 0 15792 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_133
timestamp 1663859327
transform 1 0 16240 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_139
timestamp 1663859327
transform 1 0 16912 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_147
timestamp 1663859327
transform 1 0 17808 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_155
timestamp 1663859327
transform 1 0 18704 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_159
timestamp 1663859327
transform 1 0 19152 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_163
timestamp 1663859327
transform 1 0 19600 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_167
timestamp 1663859327
transform 1 0 20048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_171
timestamp 1663859327
transform 1 0 20496 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_173
timestamp 1663859327
transform 1 0 20720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1663859327
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1663859327
transform 1 0 21392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_182
timestamp 1663859327
transform 1 0 21728 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_186
timestamp 1663859327
transform 1 0 22176 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_218
timestamp 1663859327
transform 1 0 25760 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_234
timestamp 1663859327
transform 1 0 27552 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_242
timestamp 1663859327
transform 1 0 28448 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_246
timestamp 1663859327
transform 1 0 28896 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1663859327
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1663859327
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1663859327
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1663859327
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1663859327
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1663859327
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_392
timestamp 1663859327
transform 1 0 45248 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_408
timestamp 1663859327
transform 1 0 47040 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_412
timestamp 1663859327
transform 1 0 47488 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_414
timestamp 1663859327
transform 1 0 47712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1663859327
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1663859327
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_7
timestamp 1663859327
transform 1 0 2128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_73
timestamp 1663859327
transform 1 0 9520 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_107
timestamp 1663859327
transform 1 0 13328 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_111
timestamp 1663859327
transform 1 0 13776 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_115
timestamp 1663859327
transform 1 0 14224 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_119
timestamp 1663859327
transform 1 0 14672 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_123
timestamp 1663859327
transform 1 0 15120 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_127
timestamp 1663859327
transform 1 0 15568 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_133
timestamp 1663859327
transform 1 0 16240 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1663859327
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1663859327
transform 1 0 17472 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_153
timestamp 1663859327
transform 1 0 18480 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_161
timestamp 1663859327
transform 1 0 19376 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_167
timestamp 1663859327
transform 1 0 20048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_171
timestamp 1663859327
transform 1 0 20496 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_175
timestamp 1663859327
transform 1 0 20944 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_179
timestamp 1663859327
transform 1 0 21392 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_183
timestamp 1663859327
transform 1 0 21840 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_187
timestamp 1663859327
transform 1 0 22288 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_191
timestamp 1663859327
transform 1 0 22736 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_195
timestamp 1663859327
transform 1 0 23184 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_211
timestamp 1663859327
transform 1 0 24976 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1663859327
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1663859327
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1663859327
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1663859327
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1663859327
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1663859327
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_357
timestamp 1663859327
transform 1 0 41328 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_389
timestamp 1663859327
transform 1 0 44912 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_405
timestamp 1663859327
transform 1 0 46704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_413
timestamp 1663859327
transform 1 0 47600 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_417
timestamp 1663859327
transform 1 0 48048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_419
timestamp 1663859327
transform 1 0 48272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_2
timestamp 1663859327
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1663859327
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_37
timestamp 1663859327
transform 1 0 5488 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_69
timestamp 1663859327
transform 1 0 9072 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_77
timestamp 1663859327
transform 1 0 9968 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_81
timestamp 1663859327
transform 1 0 10416 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_84
timestamp 1663859327
transform 1 0 10752 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_88
timestamp 1663859327
transform 1 0 11200 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_92
timestamp 1663859327
transform 1 0 11648 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_94
timestamp 1663859327
transform 1 0 11872 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_97
timestamp 1663859327
transform 1 0 12208 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_101
timestamp 1663859327
transform 1 0 12656 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1663859327
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_108
timestamp 1663859327
transform 1 0 13440 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_110
timestamp 1663859327
transform 1 0 13664 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_113
timestamp 1663859327
transform 1 0 14000 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_117
timestamp 1663859327
transform 1 0 14448 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_123
timestamp 1663859327
transform 1 0 15120 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_154
timestamp 1663859327
transform 1 0 18592 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_164
timestamp 1663859327
transform 1 0 19712 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_172
timestamp 1663859327
transform 1 0 20608 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1663859327
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1663859327
transform 1 0 21392 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_182
timestamp 1663859327
transform 1 0 21728 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_186
timestamp 1663859327
transform 1 0 22176 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_190
timestamp 1663859327
transform 1 0 22624 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_194
timestamp 1663859327
transform 1 0 23072 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_198
timestamp 1663859327
transform 1 0 23520 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_202
timestamp 1663859327
transform 1 0 23968 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_206
timestamp 1663859327
transform 1 0 24416 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_238
timestamp 1663859327
transform 1 0 28000 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_246
timestamp 1663859327
transform 1 0 28896 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1663859327
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1663859327
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1663859327
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1663859327
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1663859327
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1663859327
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1663859327
transform 1 0 45248 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_408
timestamp 1663859327
transform 1 0 47040 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_412
timestamp 1663859327
transform 1 0 47488 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_414
timestamp 1663859327
transform 1 0 47712 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_419
timestamp 1663859327
transform 1 0 48272 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1663859327
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_7
timestamp 1663859327
transform 1 0 2128 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_73
timestamp 1663859327
transform 1 0 9520 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_79
timestamp 1663859327
transform 1 0 10192 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_83
timestamp 1663859327
transform 1 0 10640 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_87
timestamp 1663859327
transform 1 0 11088 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_91
timestamp 1663859327
transform 1 0 11536 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_95
timestamp 1663859327
transform 1 0 11984 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_99
timestamp 1663859327
transform 1 0 12432 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_103
timestamp 1663859327
transform 1 0 12880 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_134
timestamp 1663859327
transform 1 0 16352 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1663859327
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1663859327
transform 1 0 17472 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_153
timestamp 1663859327
transform 1 0 18480 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_163
timestamp 1663859327
transform 1 0 19600 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_172
timestamp 1663859327
transform 1 0 20608 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_180
timestamp 1663859327
transform 1 0 21504 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_186
timestamp 1663859327
transform 1 0 22176 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_190
timestamp 1663859327
transform 1 0 22624 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_194
timestamp 1663859327
transform 1 0 23072 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_198
timestamp 1663859327
transform 1 0 23520 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_202
timestamp 1663859327
transform 1 0 23968 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_206
timestamp 1663859327
transform 1 0 24416 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_210
timestamp 1663859327
transform 1 0 24864 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1663859327
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1663859327
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1663859327
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1663859327
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1663859327
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1663859327
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1663859327
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_357
timestamp 1663859327
transform 1 0 41328 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_389
timestamp 1663859327
transform 1 0 44912 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_405
timestamp 1663859327
transform 1 0 46704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_413
timestamp 1663859327
transform 1 0 47600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_417
timestamp 1663859327
transform 1 0 48048 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_419
timestamp 1663859327
transform 1 0 48272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1663859327
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1663859327
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_37
timestamp 1663859327
transform 1 0 5488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_53
timestamp 1663859327
transform 1 0 7280 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_63
timestamp 1663859327
transform 1 0 8400 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_67
timestamp 1663859327
transform 1 0 8848 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_71
timestamp 1663859327
transform 1 0 9296 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_75
timestamp 1663859327
transform 1 0 9744 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_79
timestamp 1663859327
transform 1 0 10192 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_83
timestamp 1663859327
transform 1 0 10640 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_87
timestamp 1663859327
transform 1 0 11088 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_91
timestamp 1663859327
transform 1 0 11536 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_97
timestamp 1663859327
transform 1 0 12208 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1663859327
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_108
timestamp 1663859327
transform 1 0 13440 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_111
timestamp 1663859327
transform 1 0 13776 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_121
timestamp 1663859327
transform 1 0 14896 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_131
timestamp 1663859327
transform 1 0 16016 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_162
timestamp 1663859327
transform 1 0 19488 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_172
timestamp 1663859327
transform 1 0 20608 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1663859327
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1663859327
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_186
timestamp 1663859327
transform 1 0 22176 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_192
timestamp 1663859327
transform 1 0 22848 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_196
timestamp 1663859327
transform 1 0 23296 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_200
timestamp 1663859327
transform 1 0 23744 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_204
timestamp 1663859327
transform 1 0 24192 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_208
timestamp 1663859327
transform 1 0 24640 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_212
timestamp 1663859327
transform 1 0 25088 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_216
timestamp 1663859327
transform 1 0 25536 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_220
timestamp 1663859327
transform 1 0 25984 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_224
timestamp 1663859327
transform 1 0 26432 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_240
timestamp 1663859327
transform 1 0 28224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1663859327
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1663859327
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1663859327
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1663859327
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1663859327
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1663859327
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1663859327
transform 1 0 45248 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_408
timestamp 1663859327
transform 1 0 47040 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_416
timestamp 1663859327
transform 1 0 47936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_2
timestamp 1663859327
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_34
timestamp 1663859327
transform 1 0 5152 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_50
timestamp 1663859327
transform 1 0 6944 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_54
timestamp 1663859327
transform 1 0 7392 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_58
timestamp 1663859327
transform 1 0 7840 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_62
timestamp 1663859327
transform 1 0 8288 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_66
timestamp 1663859327
transform 1 0 8736 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1663859327
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_73
timestamp 1663859327
transform 1 0 9520 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_77
timestamp 1663859327
transform 1 0 9968 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_81
timestamp 1663859327
transform 1 0 10416 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_85
timestamp 1663859327
transform 1 0 10864 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_91
timestamp 1663859327
transform 1 0 11536 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_123
timestamp 1663859327
transform 1 0 15120 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_131
timestamp 1663859327
transform 1 0 16016 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1663859327
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_144
timestamp 1663859327
transform 1 0 17472 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_174
timestamp 1663859327
transform 1 0 20832 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_184
timestamp 1663859327
transform 1 0 21952 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_193
timestamp 1663859327
transform 1 0 22960 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_199
timestamp 1663859327
transform 1 0 23632 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_205
timestamp 1663859327
transform 1 0 24304 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_209
timestamp 1663859327
transform 1 0 24752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1663859327
transform 1 0 25424 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_218
timestamp 1663859327
transform 1 0 25760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_222
timestamp 1663859327
transform 1 0 26208 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_226
timestamp 1663859327
transform 1 0 26656 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_230
timestamp 1663859327
transform 1 0 27104 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_234
timestamp 1663859327
transform 1 0 27552 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_266
timestamp 1663859327
transform 1 0 31136 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_282
timestamp 1663859327
transform 1 0 32928 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1663859327
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1663859327
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1663859327
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1663859327
transform 1 0 41328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_389
timestamp 1663859327
transform 1 0 44912 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_405
timestamp 1663859327
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_413
timestamp 1663859327
transform 1 0 47600 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_419
timestamp 1663859327
transform 1 0 48272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1663859327
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1663859327
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_37
timestamp 1663859327
transform 1 0 5488 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_41
timestamp 1663859327
transform 1 0 5936 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_43
timestamp 1663859327
transform 1 0 6160 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_46
timestamp 1663859327
transform 1 0 6496 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_50
timestamp 1663859327
transform 1 0 6944 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_54
timestamp 1663859327
transform 1 0 7392 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_58
timestamp 1663859327
transform 1 0 7840 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_62
timestamp 1663859327
transform 1 0 8288 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_66
timestamp 1663859327
transform 1 0 8736 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_70
timestamp 1663859327
transform 1 0 9184 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_74
timestamp 1663859327
transform 1 0 9632 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1663859327
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_108
timestamp 1663859327
transform 1 0 13440 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_113
timestamp 1663859327
transform 1 0 14000 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_123
timestamp 1663859327
transform 1 0 15120 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_133
timestamp 1663859327
transform 1 0 16240 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_164
timestamp 1663859327
transform 1 0 19712 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_174
timestamp 1663859327
transform 1 0 20832 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1663859327
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1663859327
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_188
timestamp 1663859327
transform 1 0 22400 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_197
timestamp 1663859327
transform 1 0 23408 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_205
timestamp 1663859327
transform 1 0 24304 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_211
timestamp 1663859327
transform 1 0 24976 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_215
timestamp 1663859327
transform 1 0 25424 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_217
timestamp 1663859327
transform 1 0 25648 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_220
timestamp 1663859327
transform 1 0 25984 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_224
timestamp 1663859327
transform 1 0 26432 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_228
timestamp 1663859327
transform 1 0 26880 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_232
timestamp 1663859327
transform 1 0 27328 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_236
timestamp 1663859327
transform 1 0 27776 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_240
timestamp 1663859327
transform 1 0 28224 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1663859327
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1663859327
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1663859327
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1663859327
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1663859327
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1663859327
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_392
timestamp 1663859327
transform 1 0 45248 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_408
timestamp 1663859327
transform 1 0 47040 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_416
timestamp 1663859327
transform 1 0 47936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_2
timestamp 1663859327
transform 1 0 1568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_36
timestamp 1663859327
transform 1 0 5376 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_40
timestamp 1663859327
transform 1 0 5824 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_44
timestamp 1663859327
transform 1 0 6272 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_48
timestamp 1663859327
transform 1 0 6720 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_52
timestamp 1663859327
transform 1 0 7168 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_56
timestamp 1663859327
transform 1 0 7616 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_60
timestamp 1663859327
transform 1 0 8064 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_64
timestamp 1663859327
transform 1 0 8512 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1663859327
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_73
timestamp 1663859327
transform 1 0 9520 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_76
timestamp 1663859327
transform 1 0 9856 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_82
timestamp 1663859327
transform 1 0 10528 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_92
timestamp 1663859327
transform 1 0 11648 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_124
timestamp 1663859327
transform 1 0 15232 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_128
timestamp 1663859327
transform 1 0 15680 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1663859327
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1663859327
transform 1 0 17472 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_174
timestamp 1663859327
transform 1 0 20832 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_205
timestamp 1663859327
transform 1 0 24304 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_211
timestamp 1663859327
transform 1 0 24976 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1663859327
transform 1 0 25424 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_220
timestamp 1663859327
transform 1 0 25984 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_224
timestamp 1663859327
transform 1 0 26432 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_228
timestamp 1663859327
transform 1 0 26880 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_232
timestamp 1663859327
transform 1 0 27328 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_236
timestamp 1663859327
transform 1 0 27776 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_240
timestamp 1663859327
transform 1 0 28224 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_244
timestamp 1663859327
transform 1 0 28672 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_248
timestamp 1663859327
transform 1 0 29120 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_252
timestamp 1663859327
transform 1 0 29568 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1663859327
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1663859327
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1663859327
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_357
timestamp 1663859327
transform 1 0 41328 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_389
timestamp 1663859327
transform 1 0 44912 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_405
timestamp 1663859327
transform 1 0 46704 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_413
timestamp 1663859327
transform 1 0 47600 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_417
timestamp 1663859327
transform 1 0 48048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_419
timestamp 1663859327
transform 1 0 48272 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_2
timestamp 1663859327
transform 1 0 1568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_7
timestamp 1663859327
transform 1 0 2128 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_23
timestamp 1663859327
transform 1 0 3920 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_27
timestamp 1663859327
transform 1 0 4368 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_30
timestamp 1663859327
transform 1 0 4704 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1663859327
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_37
timestamp 1663859327
transform 1 0 5488 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_40
timestamp 1663859327
transform 1 0 5824 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_44
timestamp 1663859327
transform 1 0 6272 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_48
timestamp 1663859327
transform 1 0 6720 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_52
timestamp 1663859327
transform 1 0 7168 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_56
timestamp 1663859327
transform 1 0 7616 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_62
timestamp 1663859327
transform 1 0 8288 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_68
timestamp 1663859327
transform 1 0 8960 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_74
timestamp 1663859327
transform 1 0 9632 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1663859327
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_108
timestamp 1663859327
transform 1 0 13440 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_110
timestamp 1663859327
transform 1 0 13664 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_121
timestamp 1663859327
transform 1 0 14896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_133
timestamp 1663859327
transform 1 0 16240 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_164
timestamp 1663859327
transform 1 0 19712 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1663859327
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_179
timestamp 1663859327
transform 1 0 21392 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_209
timestamp 1663859327
transform 1 0 24752 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_218
timestamp 1663859327
transform 1 0 25760 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_226
timestamp 1663859327
transform 1 0 26656 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_232
timestamp 1663859327
transform 1 0 27328 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_236
timestamp 1663859327
transform 1 0 27776 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_240
timestamp 1663859327
transform 1 0 28224 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_244
timestamp 1663859327
transform 1 0 28672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_250
timestamp 1663859327
transform 1 0 29344 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_253
timestamp 1663859327
transform 1 0 29680 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_257
timestamp 1663859327
transform 1 0 30128 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_261
timestamp 1663859327
transform 1 0 30576 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_293
timestamp 1663859327
transform 1 0 34160 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_309
timestamp 1663859327
transform 1 0 35952 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_317
timestamp 1663859327
transform 1 0 36848 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1663859327
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1663859327
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1663859327
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_392
timestamp 1663859327
transform 1 0 45248 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_408
timestamp 1663859327
transform 1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_416
timestamp 1663859327
transform 1 0 47936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_2
timestamp 1663859327
transform 1 0 1568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_10
timestamp 1663859327
transform 1 0 2464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_16
timestamp 1663859327
transform 1 0 3136 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_20
timestamp 1663859327
transform 1 0 3584 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_24
timestamp 1663859327
transform 1 0 4032 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_28
timestamp 1663859327
transform 1 0 4480 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_32
timestamp 1663859327
transform 1 0 4928 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_36
timestamp 1663859327
transform 1 0 5376 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_40
timestamp 1663859327
transform 1 0 5824 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_44
timestamp 1663859327
transform 1 0 6272 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_50
timestamp 1663859327
transform 1 0 6944 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_56
timestamp 1663859327
transform 1 0 7616 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_62
timestamp 1663859327
transform 1 0 8288 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1663859327
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_73
timestamp 1663859327
transform 1 0 9520 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_79
timestamp 1663859327
transform 1 0 10192 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_110
timestamp 1663859327
transform 1 0 13664 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1663859327
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1663859327
transform 1 0 17472 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_174
timestamp 1663859327
transform 1 0 20832 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_205
timestamp 1663859327
transform 1 0 24304 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1663859327
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_215
timestamp 1663859327
transform 1 0 25424 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_224
timestamp 1663859327
transform 1 0 26432 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_232
timestamp 1663859327
transform 1 0 27328 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_238
timestamp 1663859327
transform 1 0 28000 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_244
timestamp 1663859327
transform 1 0 28672 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_248
timestamp 1663859327
transform 1 0 29120 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_252
timestamp 1663859327
transform 1 0 29568 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_256
timestamp 1663859327
transform 1 0 30016 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_260
timestamp 1663859327
transform 1 0 30464 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_264
timestamp 1663859327
transform 1 0 30912 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_268
timestamp 1663859327
transform 1 0 31360 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_272
timestamp 1663859327
transform 1 0 31808 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_280
timestamp 1663859327
transform 1 0 32704 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1663859327
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1663859327
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1663859327
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1663859327
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1663859327
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1663859327
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1663859327
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1663859327
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1663859327
transform 1 0 48272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1663859327
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_17
timestamp 1663859327
transform 1 0 3248 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_19
timestamp 1663859327
transform 1 0 3472 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_22
timestamp 1663859327
transform 1 0 3808 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_26
timestamp 1663859327
transform 1 0 4256 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_30
timestamp 1663859327
transform 1 0 4704 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1663859327
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_37
timestamp 1663859327
transform 1 0 5488 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_43
timestamp 1663859327
transform 1 0 6160 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_74
timestamp 1663859327
transform 1 0 9632 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1663859327
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_108
timestamp 1663859327
transform 1 0 13440 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_118
timestamp 1663859327
transform 1 0 14560 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_134
timestamp 1663859327
transform 1 0 16352 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_165
timestamp 1663859327
transform 1 0 19824 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1663859327
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_179
timestamp 1663859327
transform 1 0 21392 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_209
timestamp 1663859327
transform 1 0 24752 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_219
timestamp 1663859327
transform 1 0 25872 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_229
timestamp 1663859327
transform 1 0 26992 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_237
timestamp 1663859327
transform 1 0 27888 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_245
timestamp 1663859327
transform 1 0 28784 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1663859327
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1663859327
transform 1 0 29344 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_253
timestamp 1663859327
transform 1 0 29680 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_257
timestamp 1663859327
transform 1 0 30128 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_261
timestamp 1663859327
transform 1 0 30576 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_265
timestamp 1663859327
transform 1 0 31024 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_269
timestamp 1663859327
transform 1 0 31472 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_273
timestamp 1663859327
transform 1 0 31920 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_277
timestamp 1663859327
transform 1 0 32368 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_281
timestamp 1663859327
transform 1 0 32816 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_313
timestamp 1663859327
transform 1 0 36400 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_317
timestamp 1663859327
transform 1 0 36848 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1663859327
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1663859327
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1663859327
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_392
timestamp 1663859327
transform 1 0 45248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_408
timestamp 1663859327
transform 1 0 47040 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_416
timestamp 1663859327
transform 1 0 47936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1663859327
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_7
timestamp 1663859327
transform 1 0 2128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_13
timestamp 1663859327
transform 1 0 2800 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_17
timestamp 1663859327
transform 1 0 3248 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_21
timestamp 1663859327
transform 1 0 3696 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_25
timestamp 1663859327
transform 1 0 4144 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_29
timestamp 1663859327
transform 1 0 4592 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_33
timestamp 1663859327
transform 1 0 5040 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_39
timestamp 1663859327
transform 1 0 5712 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1663859327
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1663859327
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_82
timestamp 1663859327
transform 1 0 10528 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_94
timestamp 1663859327
transform 1 0 11872 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_126
timestamp 1663859327
transform 1 0 15456 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_128
timestamp 1663859327
transform 1 0 15680 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1663859327
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1663859327
transform 1 0 17472 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_154
timestamp 1663859327
transform 1 0 18592 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_170
timestamp 1663859327
transform 1 0 20384 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_202
timestamp 1663859327
transform 1 0 23968 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1663859327
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1663859327
transform 1 0 25424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_224
timestamp 1663859327
transform 1 0 26432 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_234
timestamp 1663859327
transform 1 0 27552 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_244
timestamp 1663859327
transform 1 0 28672 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_252
timestamp 1663859327
transform 1 0 29568 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_258
timestamp 1663859327
transform 1 0 30240 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_264
timestamp 1663859327
transform 1 0 30912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_268
timestamp 1663859327
transform 1 0 31360 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_272
timestamp 1663859327
transform 1 0 31808 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_276
timestamp 1663859327
transform 1 0 32256 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_280
timestamp 1663859327
transform 1 0 32704 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_286
timestamp 1663859327
transform 1 0 33376 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_289
timestamp 1663859327
transform 1 0 33712 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_297
timestamp 1663859327
transform 1 0 34608 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_300
timestamp 1663859327
transform 1 0 34944 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_332
timestamp 1663859327
transform 1 0 38528 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_348
timestamp 1663859327
transform 1 0 40320 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_352
timestamp 1663859327
transform 1 0 40768 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1663859327
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_357
timestamp 1663859327
transform 1 0 41328 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_389
timestamp 1663859327
transform 1 0 44912 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_405
timestamp 1663859327
transform 1 0 46704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_413
timestamp 1663859327
transform 1 0 47600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_417
timestamp 1663859327
transform 1 0 48048 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1663859327
transform 1 0 48272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1663859327
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_5
timestamp 1663859327
transform 1 0 1904 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_11
timestamp 1663859327
transform 1 0 2576 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_17
timestamp 1663859327
transform 1 0 3248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_19
timestamp 1663859327
transform 1 0 3472 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1663859327
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_37
timestamp 1663859327
transform 1 0 5488 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_39
timestamp 1663859327
transform 1 0 5712 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_69
timestamp 1663859327
transform 1 0 9072 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_72
timestamp 1663859327
transform 1 0 9408 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_74
timestamp 1663859327
transform 1 0 9632 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_104
timestamp 1663859327
transform 1 0 12992 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_107
timestamp 1663859327
transform 1 0 13328 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_138
timestamp 1663859327
transform 1 0 16800 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_142
timestamp 1663859327
transform 1 0 17248 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_173
timestamp 1663859327
transform 1 0 20720 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_177
timestamp 1663859327
transform 1 0 21168 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_208
timestamp 1663859327
transform 1 0 24640 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_212
timestamp 1663859327
transform 1 0 25088 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_242
timestamp 1663859327
transform 1 0 28448 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_244
timestamp 1663859327
transform 1 0 28672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1663859327
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_256
timestamp 1663859327
transform 1 0 30016 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_262
timestamp 1663859327
transform 1 0 30688 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_264
timestamp 1663859327
transform 1 0 30912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_271
timestamp 1663859327
transform 1 0 31696 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_275
timestamp 1663859327
transform 1 0 32144 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_279
timestamp 1663859327
transform 1 0 32592 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_282
timestamp 1663859327
transform 1 0 32928 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_297
timestamp 1663859327
transform 1 0 34608 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_299
timestamp 1663859327
transform 1 0 34832 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_314
timestamp 1663859327
transform 1 0 36512 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_317
timestamp 1663859327
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_329
timestamp 1663859327
transform 1 0 38192 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_337
timestamp 1663859327
transform 1 0 39088 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_341
timestamp 1663859327
transform 1 0 39536 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_347
timestamp 1663859327
transform 1 0 40208 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_349
timestamp 1663859327
transform 1 0 40432 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_352
timestamp 1663859327
transform 1 0 40768 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_360
timestamp 1663859327
transform 1 0 41664 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_364
timestamp 1663859327
transform 1 0 42112 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_368
timestamp 1663859327
transform 1 0 42560 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_384
timestamp 1663859327
transform 1 0 44352 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_387
timestamp 1663859327
transform 1 0 44688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_403
timestamp 1663859327
transform 1 0 46480 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_411
timestamp 1663859327
transform 1 0 47376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_419
timestamp 1663859327
transform 1 0 48272 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1663859327
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1663859327
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1663859327
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1663859327
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1663859327
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1663859327
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1663859327
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1663859327
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1663859327
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1663859327
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1663859327
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1663859327
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1663859327
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1663859327
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1663859327
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1663859327
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1663859327
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1663859327
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1663859327
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1663859327
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1663859327
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1663859327
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1663859327
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1663859327
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1663859327
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1663859327
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1663859327
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1663859327
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1663859327
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1663859327
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1663859327
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1663859327
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1663859327
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1663859327
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1663859327
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1663859327
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1663859327
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1663859327
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1663859327
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1663859327
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1663859327
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1663859327
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1663859327
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1663859327
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1663859327
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1663859327
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1663859327
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1663859327
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1663859327
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1663859327
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1663859327
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1663859327
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1663859327
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1663859327
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1663859327
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1663859327
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1663859327
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1663859327
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1663859327
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1663859327
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1663859327
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1663859327
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1663859327
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1663859327
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1663859327
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1663859327
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1663859327
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1663859327
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1663859327
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1663859327
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1663859327
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1663859327
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1663859327
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1663859327
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1663859327
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1663859327
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1663859327
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1663859327
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1663859327
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1663859327
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1663859327
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1663859327
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1663859327
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1663859327
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1663859327
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1663859327
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1663859327
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1663859327
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1663859327
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1663859327
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1663859327
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1663859327
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1663859327
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1663859327
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1663859327
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1663859327
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1663859327
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1663859327
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1663859327
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1663859327
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1663859327
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1663859327
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1663859327
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1663859327
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1663859327
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1663859327
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1663859327
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1663859327
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1663859327
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1663859327
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1663859327
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1663859327
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1663859327
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1663859327
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1663859327
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1663859327
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1663859327
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1663859327
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1663859327
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1663859327
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1663859327
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1663859327
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1663859327
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1663859327
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1663859327
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1663859327
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1663859327
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1663859327
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1663859327
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1663859327
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1663859327
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1663859327
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1663859327
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1663859327
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1663859327
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1663859327
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1663859327
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1663859327
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1663859327
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1663859327
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1663859327
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1663859327
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1663859327
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1663859327
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1663859327
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1663859327
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1663859327
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1663859327
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1663859327
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1663859327
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1663859327
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1663859327
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1663859327
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1663859327
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1663859327
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1663859327
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1663859327
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1663859327
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1663859327
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1663859327
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1663859327
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1663859327
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1663859327
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1663859327
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1663859327
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1663859327
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1663859327
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1663859327
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1663859327
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1663859327
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1663859327
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1663859327
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1663859327
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1663859327
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1663859327
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1663859327
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1663859327
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1663859327
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1663859327
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1663859327
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1663859327
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1663859327
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1663859327
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1663859327
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1663859327
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1663859327
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1663859327
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1663859327
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1663859327
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1663859327
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1663859327
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1663859327
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1663859327
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1663859327
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1663859327
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1663859327
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1663859327
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1663859327
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1663859327
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1663859327
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1663859327
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1663859327
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1663859327
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1663859327
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1663859327
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1663859327
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1663859327
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1663859327
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1663859327
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1663859327
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1663859327
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1663859327
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1663859327
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1663859327
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1663859327
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1663859327
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1663859327
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1663859327
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1663859327
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1663859327
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1663859327
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1663859327
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1663859327
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1663859327
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1663859327
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1663859327
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1663859327
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1663859327
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1663859327
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1663859327
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1663859327
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1663859327
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1663859327
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1663859327
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1663859327
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1663859327
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1663859327
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1663859327
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1663859327
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1663859327
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1663859327
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1663859327
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1663859327
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1663859327
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1663859327
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1663859327
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1663859327
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1663859327
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1663859327
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1663859327
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1663859327
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1663859327
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1663859327
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1663859327
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1663859327
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1663859327
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1663859327
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1663859327
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1663859327
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1663859327
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1663859327
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1663859327
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1663859327
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1663859327
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1663859327
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1663859327
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1663859327
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1663859327
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1663859327
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1663859327
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1663859327
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1663859327
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1663859327
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1663859327
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1663859327
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1663859327
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1663859327
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1663859327
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1663859327
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1663859327
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1663859327
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1663859327
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1663859327
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1663859327
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1663859327
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1663859327
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1663859327
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1663859327
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1663859327
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1663859327
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1663859327
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1663859327
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1663859327
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1663859327
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1663859327
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1663859327
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1663859327
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1663859327
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1663859327
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1663859327
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1663859327
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1663859327
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1663859327
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1663859327
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1663859327
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1663859327
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1663859327
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1663859327
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1663859327
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1663859327
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1663859327
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1663859327
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1663859327
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1663859327
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1663859327
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1663859327
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1663859327
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1663859327
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1663859327
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1663859327
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1663859327
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1663859327
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1663859327
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1663859327
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1663859327
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1663859327
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1663859327
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1663859327
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1663859327
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1663859327
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1663859327
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1663859327
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1663859327
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1663859327
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1663859327
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1663859327
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1663859327
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1663859327
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1663859327
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1663859327
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1663859327
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1663859327
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1663859327
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1663859327
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1663859327
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1663859327
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1663859327
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1663859327
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1663859327
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1663859327
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1663859327
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1663859327
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1663859327
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1663859327
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1663859327
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1663859327
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1663859327
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1663859327
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1663859327
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1663859327
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1663859327
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1663859327
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1663859327
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1663859327
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1663859327
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1663859327
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1663859327
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1663859327
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1663859327
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1663859327
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1663859327
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1663859327
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1663859327
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1663859327
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1663859327
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1663859327
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1663859327
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1663859327
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1663859327
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1663859327
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1663859327
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1663859327
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1663859327
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1663859327
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1663859327
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1663859327
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1663859327
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1663859327
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1663859327
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1663859327
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1663859327
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1663859327
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1663859327
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1663859327
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1663859327
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1663859327
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1663859327
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1663859327
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1663859327
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1663859327
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1663859327
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1663859327
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1663859327
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1663859327
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1663859327
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1663859327
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1663859327
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1663859327
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1663859327
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1663859327
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1663859327
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1663859327
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1663859327
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1663859327
transform 1 0 17024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1663859327
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1663859327
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1663859327
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1663859327
transform 1 0 32704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1663859327
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1663859327
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1663859327
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _050_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 9184 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _051_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 24304 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _052_
timestamp 1663859327
transform 1 0 7840 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _053_
timestamp 1663859327
transform -1 0 10528 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _054_
timestamp 1663859327
transform -1 0 25984 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _055_
timestamp 1663859327
transform 1 0 23184 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _056_
timestamp 1663859327
transform 1 0 5264 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _057_
timestamp 1663859327
transform 1 0 20832 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _058_
timestamp 1663859327
transform -1 0 13104 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _059_
timestamp 1663859327
transform 1 0 15792 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _060_
timestamp 1663859327
transform 1 0 28224 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _061_
timestamp 1663859327
transform -1 0 22176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _062_
timestamp 1663859327
transform -1 0 24304 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _063_
timestamp 1663859327
transform -1 0 24976 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _064_
timestamp 1663859327
transform 1 0 19600 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _065_
timestamp 1663859327
transform -1 0 27328 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _066_
timestamp 1663859327
transform -1 0 30240 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _067_
timestamp 1663859327
transform -1 0 16912 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _068_
timestamp 1663859327
transform -1 0 11536 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _069_
timestamp 1663859327
transform 1 0 5712 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _070_
timestamp 1663859327
transform 1 0 7840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _071_
timestamp 1663859327
transform -1 0 24976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _072_
timestamp 1663859327
transform -1 0 18704 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _073_
timestamp 1663859327
transform 1 0 27216 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _074_
timestamp 1663859327
transform -1 0 22176 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _075_
timestamp 1663859327
transform 1 0 7168 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _076_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 16576 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _077_
timestamp 1663859327
transform -1 0 26656 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _078_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 8512 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _079_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 25760 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _080_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 17584 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _081_
timestamp 1663859327
transform 1 0 27552 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _082_
timestamp 1663859327
transform -1 0 20608 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _083_
timestamp 1663859327
transform 1 0 16464 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _084_
timestamp 1663859327
transform 1 0 8512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _085_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 13552 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _086_
timestamp 1663859327
transform -1 0 15120 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _087_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 26096 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _088_
timestamp 1663859327
transform -1 0 17808 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _089_
timestamp 1663859327
transform -1 0 10528 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _090_
timestamp 1663859327
transform -1 0 19376 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _091_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 15120 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _092_
timestamp 1663859327
transform -1 0 18480 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _093_
timestamp 1663859327
transform 1 0 17584 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _094_
timestamp 1663859327
transform -1 0 20832 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _095_
timestamp 1663859327
transform -1 0 23408 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _096_
timestamp 1663859327
transform 1 0 18704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _097_
timestamp 1663859327
transform 1 0 25536 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _098_
timestamp 1663859327
transform 1 0 14000 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _099_
timestamp 1663859327
transform -1 0 16016 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _100_
timestamp 1663859327
transform 1 0 28112 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _101_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 16240 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _102_
timestamp 1663859327
transform 1 0 26656 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _103_
timestamp 1663859327
transform 1 0 16240 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _104_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 17136 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _105_
timestamp 1663859327
transform -1 0 10192 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _106_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 11872 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _107_
timestamp 1663859327
transform -1 0 30016 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _108_
timestamp 1663859327
transform 1 0 21504 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _109_
timestamp 1663859327
transform -1 0 21056 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _110_
timestamp 1663859327
transform -1 0 26432 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _111_
timestamp 1663859327
transform -1 0 21952 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _112_
timestamp 1663859327
transform 1 0 24976 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _113_
timestamp 1663859327
transform 1 0 26656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _114_
timestamp 1663859327
transform 1 0 13776 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _115_
timestamp 1663859327
transform -1 0 25088 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _116_
timestamp 1663859327
transform -1 0 16016 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _117_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 21056 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _118_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 16352 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _119_
timestamp 1663859327
transform -1 0 22960 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _120_
timestamp 1663859327
transform 1 0 18816 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _121_
timestamp 1663859327
transform -1 0 20608 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _122_
timestamp 1663859327
transform 1 0 27776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _123_
timestamp 1663859327
transform -1 0 15120 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _124_
timestamp 1663859327
transform -1 0 29568 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _125_
timestamp 1663859327
transform 1 0 15792 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1663859327
transform 1 0 19936 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1663859327
transform 1 0 30464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _128_
timestamp 1663859327
transform 1 0 24192 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _129_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 20608 0 -1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _130_
timestamp 1663859327
transform -1 0 20720 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _131_
timestamp 1663859327
transform -1 0 16800 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _132_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 16576 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _133_
timestamp 1663859327
transform 1 0 17584 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _134_
timestamp 1663859327
transform -1 0 19712 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _135_
timestamp 1663859327
transform -1 0 24304 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _136_
timestamp 1663859327
transform 1 0 16240 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _137_
timestamp 1663859327
transform -1 0 24752 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _138_
timestamp 1663859327
transform 1 0 21504 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _139_
timestamp 1663859327
transform -1 0 17136 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _140_
timestamp 1663859327
transform -1 0 20832 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _141_
timestamp 1663859327
transform -1 0 20832 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _142_
timestamp 1663859327
transform -1 0 28448 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _143_
timestamp 1663859327
transform 1 0 9744 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _144_
timestamp 1663859327
transform -1 0 13104 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _145_
timestamp 1663859327
transform 1 0 15344 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _146_
timestamp 1663859327
transform 1 0 6384 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _147_
timestamp 1663859327
transform 1 0 13104 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _148_
timestamp 1663859327
transform 1 0 9856 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _149_
timestamp 1663859327
transform -1 0 19712 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _150_
timestamp 1663859327
transform 1 0 10416 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _151_
timestamp 1663859327
transform 1 0 21280 0 1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _152_
timestamp 1663859327
transform -1 0 13104 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _153_
timestamp 1663859327
transform -1 0 9072 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _154_
timestamp 1663859327
transform 1 0 5936 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _155_
timestamp 1663859327
transform -1 0 24304 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _156_
timestamp 1663859327
transform -1 0 15232 0 -1 42336
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _157_
timestamp 1663859327
transform -1 0 15120 0 -1 40768
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _158_
timestamp 1663859327
transform -1 0 15456 0 -1 45472
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input1 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 10752 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1663859327
transform -1 0 31696 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output3 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 5152 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output4
timestamp 1663859327
transform 1 0 18816 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output5
timestamp 1663859327
transform 1 0 34944 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output6
timestamp 1663859327
transform -1 0 3248 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output7
timestamp 1663859327
transform -1 0 3248 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output8
timestamp 1663859327
transform -1 0 3248 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output9
timestamp 1663859327
transform 1 0 42784 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output10
timestamp 1663859327
transform 1 0 33040 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_11 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 2128 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_12
timestamp 1663859327
transform -1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_13
timestamp 1663859327
transform 1 0 47824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_14
timestamp 1663859327
transform -1 0 38192 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_15
timestamp 1663859327
transform -1 0 2576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_16
timestamp 1663859327
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_17
timestamp 1663859327
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_18
timestamp 1663859327
transform -1 0 2128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_19
timestamp 1663859327
transform -1 0 2128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_20
timestamp 1663859327
transform 1 0 47824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_21
timestamp 1663859327
transform -1 0 2128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_22
timestamp 1663859327
transform -1 0 2128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_23
timestamp 1663859327
transform 1 0 47824 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_24
timestamp 1663859327
transform 1 0 47824 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_25
timestamp 1663859327
transform -1 0 42896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_26
timestamp 1663859327
transform 1 0 47824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_27
timestamp 1663859327
transform -1 0 2128 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_28
timestamp 1663859327
transform -1 0 2128 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_29
timestamp 1663859327
transform -1 0 26768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_30
timestamp 1663859327
transform -1 0 2800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_31
timestamp 1663859327
transform -1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_32
timestamp 1663859327
transform 1 0 47824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_33
timestamp 1663859327
transform -1 0 3248 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_34
timestamp 1663859327
transform -1 0 2128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_35
timestamp 1663859327
transform -1 0 9968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_36
timestamp 1663859327
transform -1 0 18032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_37
timestamp 1663859327
transform -1 0 2128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_38
timestamp 1663859327
transform 1 0 47824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_39
timestamp 1663859327
transform -1 0 29568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_40
timestamp 1663859327
transform -1 0 40208 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_41
timestamp 1663859327
transform -1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_42
timestamp 1663859327
transform -1 0 30688 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_43
timestamp 1663859327
transform -1 0 41328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_44
timestamp 1663859327
transform -1 0 2128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_45
timestamp 1663859327
transform -1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_46
timestamp 1663859327
transform -1 0 2128 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_47
timestamp 1663859327
transform 1 0 47824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_48
timestamp 1663859327
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_49
timestamp 1663859327
transform 1 0 47824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_50
timestamp 1663859327
transform -1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_51
timestamp 1663859327
transform -1 0 2128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_52
timestamp 1663859327
transform 1 0 47824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_53
timestamp 1663859327
transform -1 0 2128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_54
timestamp 1663859327
transform -1 0 2128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_55
timestamp 1663859327
transform 1 0 47824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_56
timestamp 1663859327
transform -1 0 44240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_57
timestamp 1663859327
transform -1 0 2128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_58
timestamp 1663859327
transform 1 0 47824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_59
timestamp 1663859327
transform -1 0 22848 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_60
timestamp 1663859327
transform 1 0 11760 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_61
timestamp 1663859327
transform 1 0 13552 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_62
timestamp 1663859327
transform -1 0 14672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_63
timestamp 1663859327
transform 1 0 47824 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_64
timestamp 1663859327
transform 1 0 47824 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_65
timestamp 1663859327
transform 1 0 47824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_66
timestamp 1663859327
transform -1 0 3920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_67
timestamp 1663859327
transform -1 0 46256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_68
timestamp 1663859327
transform 1 0 47824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_69
timestamp 1663859327
transform -1 0 2128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_70
timestamp 1663859327
transform -1 0 2128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_71
timestamp 1663859327
transform -1 0 21728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_72
timestamp 1663859327
transform 1 0 47824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_73
timestamp 1663859327
transform 1 0 47824 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_74
timestamp 1663859327
transform -1 0 2128 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_75
timestamp 1663859327
transform 1 0 47152 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_76
timestamp 1663859327
transform -1 0 2800 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_77
timestamp 1663859327
transform 1 0 6496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_78
timestamp 1663859327
transform -1 0 2128 0 1 32928
box -86 -86 534 870
<< labels >>
flabel metal2 s 23520 49200 23632 49800 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 49728 49200 49840 49800 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 24192 200 24304 800 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 11424 49200 11536 49800 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 49056 200 49168 800 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 49200 43008 49800 43120 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 36960 200 37072 800 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 12096 200 12208 800 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 200 47712 800 47824 0 FreeSans 448 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 18816 200 18928 800 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30912 49200 31024 49800 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 200 1344 800 1456 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 33600 200 33712 800 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal3 s 200 31584 800 31696 0 FreeSans 448 0 0 0 io_in[21]
port 13 nsew signal input
flabel metal3 s 49200 20160 49800 20272 0 FreeSans 448 0 0 0 io_in[22]
port 14 nsew signal input
flabel metal3 s 49200 46368 49800 46480 0 FreeSans 448 0 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 200 4704 800 4816 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 40992 49200 41104 49800 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 200 40320 800 40432 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 49200 14784 49800 14896 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 49200 40992 49800 41104 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 47712 200 47824 800 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 29568 200 29680 800 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 49200 4032 49800 4144 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 14784 49200 14896 49800 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 10080 200 10192 800 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 25536 49200 25648 49800 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 46368 49200 46480 49800 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 200 12096 800 12208 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 16128 49200 16240 49800 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 49200 45024 49800 45136 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 49200 25536 49800 25648 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 28896 49200 29008 49800 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 6720 200 6832 800 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 45024 49200 45136 49800 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 34272 49200 34384 49800 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 6048 49200 6160 49800 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 49200 48384 49800 48496 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 15456 200 15568 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 200 8736 800 8848 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 49200 34272 49800 34384 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 200 34944 800 35056 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 200 18816 800 18928 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 49200 11424 49800 11536 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 43680 200 43792 800 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal3 s 200 24192 800 24304 0 FreeSans 448 0 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal3 s 49200 26880 49800 26992 0 FreeSans 448 0 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 21504 49200 21616 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 12768 49200 12880 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 26880 49200 26992 49800 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 18144 49200 18256 49800 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 14112 200 14224 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal3 s 49200 12768 49800 12880 0 FreeSans 448 0 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal3 s 49200 6048 49800 6160 0 FreeSans 448 0 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 49200 32256 49800 32368 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 3360 200 3472 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 45696 200 45808 800 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 49200 9408 49800 9520 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 200 29568 800 29680 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 200 3360 800 3472 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 40320 200 40432 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 20832 200 20944 800 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 49200 16800 49800 16912 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 49200 37632 49800 37744 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 200 38304 800 38416 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 49200 2016 49800 2128 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 200 45696 800 45808 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 7392 49200 7504 49800 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 200 32928 800 33040 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 200 6720 800 6832 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 4704 200 4816 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 200 20832 800 20944 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 49200 672 49800 784 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 49200 28896 49800 29008 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 49200 18144 49800 18256 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 38304 200 38416 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 200 36960 800 37072 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 200 28224 800 28336 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 200 26208 800 26320 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 49200 21504 49800 21616 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 49200 35616 49800 35728 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 42336 200 42448 800 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal3 s 49200 39648 49800 39760 0 FreeSans 448 0 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 672 49200 784 49800 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal3 s 200 10080 800 10192 0 FreeSans 448 0 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 26208 200 26320 800 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 31584 200 31696 800 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 4032 49200 4144 49800 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 20160 49200 20272 49800 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35616 49200 35728 49800 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal3 s 200 43680 800 43792 0 FreeSans 448 0 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 200 22848 800 22960 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 1344 200 1456 800 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 43008 49200 43120 49800 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 32256 49200 32368 49800 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 22848 200 22960 800 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 48384 49200 48496 49800 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 49200 7392 49800 7504 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 200 49056 800 49168 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 200 17472 800 17584 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 8736 200 8848 800 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 17472 200 17584 800 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 200 15456 800 15568 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 49200 30912 49800 31024 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 28224 200 28336 800 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 39648 49200 39760 49800 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 37632 49200 37744 49800 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 2016 49200 2128 49800 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 9408 49200 9520 49800 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 34944 200 35056 800 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 200 14112 800 14224 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 200 42336 800 42448 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 49200 23520 49800 23632 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vccd1
rlabel metal1 24976 45472 24976 45472 0 vssd1
rlabel metal2 24472 45416 24472 45416 0 _000_
rlabel metal3 21000 39032 21000 39032 0 _001_
rlabel metal2 21784 40264 21784 40264 0 _002_
rlabel metal2 25760 43736 25760 43736 0 _003_
rlabel metal2 16296 45584 16296 45584 0 _004_
rlabel metal2 22344 42616 22344 42616 0 _005_
rlabel metal2 15512 41440 15512 41440 0 _006_
rlabel metal3 25256 43456 25256 43456 0 _007_
rlabel metal2 16520 42672 16520 42672 0 _008_
rlabel metal3 13720 44968 13720 44968 0 _009_
rlabel metal2 24696 39704 24696 39704 0 _010_
rlabel metal2 26264 45472 26264 45472 0 _011_
rlabel metal2 21784 41664 21784 41664 0 _012_
rlabel metal2 25592 43456 25592 43456 0 _013_
rlabel metal2 25144 43904 25144 43904 0 _014_
rlabel metal2 14168 43288 14168 43288 0 _015_
rlabel metal2 24584 43848 24584 43848 0 _016_
rlabel metal2 15736 39816 15736 39816 0 _017_
rlabel metal2 19992 39872 19992 39872 0 _018_
rlabel metal3 18816 38696 18816 38696 0 _019_
rlabel metal4 20328 40992 20328 40992 0 _020_
rlabel metal2 15008 37912 15008 37912 0 _021_
rlabel metal2 16744 42728 16744 42728 0 _022_
rlabel metal2 20048 38024 20048 38024 0 _023_
rlabel metal2 18424 45304 18424 45304 0 _024_
rlabel metal2 16408 45360 16408 45360 0 _025_
rlabel metal2 10640 38136 10640 38136 0 _026_
rlabel metal2 24920 40264 24920 40264 0 _027_
rlabel metal2 25312 44072 25312 44072 0 _028_
rlabel metal2 26712 43736 26712 43736 0 _029_
rlabel metal2 18704 35000 18704 35000 0 _030_
rlabel metal2 14728 36792 14728 36792 0 _031_
rlabel metal3 18312 38808 18312 38808 0 _032_
rlabel metal2 25816 40880 25816 40880 0 _033_
rlabel metal3 22512 41160 22512 41160 0 _034_
rlabel metal2 18424 39088 18424 39088 0 _035_
rlabel metal2 29400 40432 29400 40432 0 _036_
rlabel metal2 18200 44520 18200 44520 0 _037_
rlabel metal2 20720 40936 20720 40936 0 _038_
rlabel metal2 16408 41888 16408 41888 0 _039_
rlabel metal2 17752 44128 17752 44128 0 _040_
rlabel metal2 14280 42840 14280 42840 0 _041_
rlabel metal4 26824 44184 26824 44184 0 _042_
rlabel metal2 26544 42840 26544 42840 0 _043_
rlabel metal2 20888 42840 20888 42840 0 _044_
rlabel metal2 15736 42784 15736 42784 0 _045_
rlabel metal2 20104 42784 20104 42784 0 _046_
rlabel metal2 14840 39368 14840 39368 0 _047_
rlabel metal2 19992 41608 19992 41608 0 _048_
rlabel metal2 20608 41160 20608 41160 0 _049_
rlabel metal2 8736 40600 8736 40600 0 io_in[12]
rlabel metal2 31416 46032 31416 46032 0 io_in[19]
rlabel metal2 4088 47642 4088 47642 0 io_out[20]
rlabel metal2 20104 44968 20104 44968 0 io_out[21]
rlabel metal2 35728 45976 35728 45976 0 io_out[22]
rlabel metal3 1470 43736 1470 43736 0 io_out[23]
rlabel metal3 1414 22904 1414 22904 0 io_out[24]
rlabel metal2 1400 2142 1400 2142 0 io_out[25]
rlabel metal2 43064 47642 43064 47642 0 io_out[26]
rlabel metal3 33096 45976 33096 45976 0 io_out[27]
rlabel metal2 10808 41888 10808 41888 0 mod.flipflop1.d
rlabel metal2 12600 38192 12600 38192 0 mod.flipflop1.q
rlabel metal2 17752 41944 17752 41944 0 mod.flipflop10.clk
rlabel metal2 21896 39088 21896 39088 0 mod.flipflop10.d
rlabel metal2 21672 43904 21672 43904 0 mod.flipflop10.q
rlabel metal2 22456 44072 22456 44072 0 mod.flipflop11.d
rlabel metal2 24640 44408 24640 44408 0 mod.flipflop11.q
rlabel metal2 23744 42616 23744 42616 0 mod.flipflop12.d
rlabel metal2 13048 37464 13048 37464 0 mod.flipflop12.q
rlabel metal2 11032 38360 11032 38360 0 mod.flipflop13.d
rlabel metal2 24248 43512 24248 43512 0 mod.flipflop13.q
rlabel metal2 15232 39480 15232 39480 0 mod.flipflop14.d
rlabel metal2 21224 43176 21224 43176 0 mod.flipflop14.q
rlabel metal3 22232 41272 22232 41272 0 mod.flipflop15.d
rlabel metal2 16632 41384 16632 41384 0 mod.flipflop15.q
rlabel metal2 18536 42672 18536 42672 0 mod.flipflop16.d
rlabel metal2 20664 43624 20664 43624 0 mod.flipflop16.q
rlabel metal2 15624 39648 15624 39648 0 mod.flipflop17.d
rlabel metal2 19656 44968 19656 44968 0 mod.flipflop17.q
rlabel metal2 14504 44352 14504 44352 0 mod.flipflop18.d
rlabel metal2 25256 45136 25256 45136 0 mod.flipflop19.d
rlabel metal3 8680 39032 8680 39032 0 mod.flipflop2.d
rlabel metal2 16184 38808 16184 38808 0 mod.flipflop2.q
rlabel metal3 23800 45080 23800 45080 0 mod.flipflop20.d
rlabel metal3 12880 45080 12880 45080 0 mod.flipflop21.d
rlabel metal2 14280 40040 14280 40040 0 mod.flipflop22.d
rlabel metal2 18144 37464 18144 37464 0 mod.flipflop23.d
rlabel metal2 23296 40488 23296 40488 0 mod.flipflop25.d
rlabel metal2 21168 41832 21168 41832 0 mod.flipflop25.q
rlabel metal2 18760 42224 18760 42224 0 mod.flipflop26.d
rlabel metal2 16632 43064 16632 43064 0 mod.flipflop26.q
rlabel metal2 24248 46648 24248 46648 0 mod.flipflop27.d
rlabel metal2 16296 42840 16296 42840 0 mod.flipflop27.q
rlabel metal3 10640 37912 10640 37912 0 mod.flipflop28.d
rlabel metal3 27412 36792 27412 36792 0 mod.flipflop28.q
rlabel metal2 19096 37744 19096 37744 0 mod.flipflop29.d
rlabel metal2 26712 41776 26712 41776 0 mod.flipflop29.q
rlabel metal2 11256 42392 11256 42392 0 mod.flipflop3.d
rlabel metal3 13048 37464 13048 37464 0 mod.flipflop3.q
rlabel metal2 16744 46592 16744 46592 0 mod.flipflop30.q
rlabel metal2 16576 36680 16576 36680 0 mod.flipflop4.d
rlabel metal2 15848 39872 15848 39872 0 mod.flipflop4.q
rlabel metal2 20328 45752 20328 45752 0 mod.flipflop5.d
rlabel metal2 10024 46816 10024 46816 0 mod.flipflop5.q
rlabel metal2 25480 45584 25480 45584 0 mod.flipflop6.d
rlabel metal2 24920 45080 24920 45080 0 mod.flipflop6.q
rlabel metal2 19432 42700 19432 42700 0 mod.flipflop7.d
rlabel metal2 20664 40488 20664 40488 0 mod.flipflop7.q
rlabel metal2 19880 40544 19880 40544 0 mod.flipflop8.d
rlabel metal2 20552 41664 20552 41664 0 mod.flipflop8.q
rlabel metal2 24024 40768 24024 40768 0 mod.flipflop9.d
rlabel metal2 24136 41496 24136 41496 0 net1
rlabel metal2 20552 45752 20552 45752 0 net10
rlabel metal3 1302 37016 1302 37016 0 net11
rlabel metal2 31640 2030 31640 2030 0 net12
rlabel metal2 48104 7728 48104 7728 0 net13
rlabel metal2 37800 45752 37800 45752 0 net14
rlabel metal2 2184 45752 2184 45752 0 net15
rlabel metal2 9072 42168 9072 42168 0 net16
rlabel metal2 35000 2030 35000 2030 0 net17
rlabel metal3 1302 14168 1302 14168 0 net18
rlabel metal3 1302 42392 1302 42392 0 net19
rlabel metal2 25368 41552 25368 41552 0 net2
rlabel metal2 48104 23632 48104 23632 0 net20
rlabel metal3 1302 28280 1302 28280 0 net21
rlabel metal3 1302 26264 1302 26264 0 net22
rlabel metal2 48104 21840 48104 21840 0 net23
rlabel metal2 48104 35952 48104 35952 0 net24
rlabel metal2 42392 2030 42392 2030 0 net25
rlabel metal2 48104 40096 48104 40096 0 net26
rlabel metal2 1792 45304 1792 45304 0 net27
rlabel metal3 1302 10136 1302 10136 0 net28
rlabel metal2 26264 2030 26264 2030 0 net29
rlabel metal3 9296 45864 9296 45864 0 net3
rlabel metal2 56 1526 56 1526 0 net30
rlabel metal2 22904 2030 22904 2030 0 net31
rlabel metal2 48272 45752 48272 45752 0 net32
rlabel metal2 2968 46368 2968 46368 0 net33
rlabel metal3 1302 17528 1302 17528 0 net34
rlabel metal2 8792 1246 8792 1246 0 net35
rlabel metal2 17528 2030 17528 2030 0 net36
rlabel metal3 1302 15512 1302 15512 0 net37
rlabel metal2 48104 31248 48104 31248 0 net38
rlabel metal2 28280 2030 28280 2030 0 net39
rlabel metal2 18984 45360 18984 45360 0 net4
rlabel metal2 39816 45752 39816 45752 0 net40
rlabel metal2 15512 2030 15512 2030 0 net41
rlabel metal3 28672 45752 28672 45752 0 net42
rlabel metal2 40376 1302 40376 1302 0 net43
rlabel metal3 1302 6776 1302 6776 0 net44
rlabel metal2 4760 2030 4760 2030 0 net45
rlabel metal3 1302 20888 1302 20888 0 net46
rlabel metal2 48104 2016 48104 2016 0 net47
rlabel metal2 48104 29232 48104 29232 0 net48
rlabel metal3 48104 18368 48104 18368 0 net49
rlabel metal2 35112 45584 35112 45584 0 net5
rlabel metal2 38360 2030 38360 2030 0 net50
rlabel metal3 1302 8792 1302 8792 0 net51
rlabel metal2 48104 34496 48104 34496 0 net52
rlabel metal3 1302 35000 1302 35000 0 net53
rlabel metal3 1302 18872 1302 18872 0 net54
rlabel metal2 48104 11872 48104 11872 0 net55
rlabel metal2 43736 2030 43736 2030 0 net56
rlabel metal3 1302 24248 1302 24248 0 net57
rlabel metal3 48104 26880 48104 26880 0 net58
rlabel metal2 22512 39480 22512 39480 0 net59
rlabel metal2 3080 45360 3080 45360 0 net6
rlabel metal2 12040 40544 12040 40544 0 net60
rlabel metal2 18088 43792 18088 43792 0 net61
rlabel metal2 14168 2030 14168 2030 0 net62
rlabel metal3 48706 12824 48706 12824 0 net63
rlabel metal2 48104 6272 48104 6272 0 net64
rlabel metal2 48104 32480 48104 32480 0 net65
rlabel metal2 3416 2030 3416 2030 0 net66
rlabel metal2 45752 2030 45752 2030 0 net67
rlabel metal2 48104 9520 48104 9520 0 net68
rlabel metal3 1302 29624 1302 29624 0 net69
rlabel metal2 3080 23240 3080 23240 0 net7
rlabel metal3 1302 3416 1302 3416 0 net70
rlabel metal2 20888 1246 20888 1246 0 net71
rlabel metal2 48104 17136 48104 17136 0 net72
rlabel metal2 48104 37744 48104 37744 0 net73
rlabel metal3 1302 38360 1302 38360 0 net74
rlabel metal2 47432 2688 47432 2688 0 net75
rlabel metal2 2520 45528 2520 45528 0 net76
rlabel metal2 6776 43792 6776 43792 0 net77
rlabel metal3 1302 32984 1302 32984 0 net78
rlabel metal3 5096 3640 5096 3640 0 net8
rlabel metal2 42504 46200 42504 46200 0 net9
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
